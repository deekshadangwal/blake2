
module blake2 ( clk, reset_n, cs, we, address, write_data, read_data, error );
  input [7:0] address;
  input [31:0] write_data;
  output [31:0] read_data;
  input clk, reset_n, cs, we;
  output error;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, read_data_30, read_data_26,
         read_data_8, read_data_6, read_data_5, read_data_4, read_data_1,
         read_data_0, core_init, core_next, core_ready, core_digest_valid,
         ready_reg, digest_valid_reg, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N128, N129, N138, N139,
         N140, N141, N142, N143, N144, N147, N148, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N161, N162, N163, N164, N165,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237;
  wire   [1023:0] core_block;
  assign read_data[2] = 1'b0;
  assign read_data[7] = 1'b0;
  assign read_data[9] = 1'b0;
  assign read_data[10] = 1'b0;
  assign read_data[11] = 1'b0;
  assign read_data[15] = 1'b0;
  assign read_data[16] = 1'b0;
  assign read_data[23] = 1'b0;
  assign read_data[27] = 1'b0;
  assign read_data[31] = 1'b0;
  assign read_data[30] = read_data_30;
  assign read_data[24] = read_data_26;
  assign read_data[20] = read_data_26;
  assign read_data[26] = read_data_26;
  assign read_data[19] = read_data_8;
  assign read_data[18] = read_data_8;
  assign read_data[8] = read_data_8;
  assign read_data[3] = read_data_6;
  assign read_data[14] = read_data_6;
  assign read_data[22] = read_data_6;
  assign read_data[25] = read_data_6;
  assign read_data[6] = read_data_6;
  assign read_data[29] = read_data_5;
  assign read_data[21] = read_data_5;
  assign read_data[13] = read_data_5;
  assign read_data[5] = read_data_5;
  assign read_data[28] = read_data_4;
  assign read_data[12] = read_data_4;
  assign read_data[4] = read_data_4;
  assign read_data[1] = read_data_1;
  assign read_data[0] = read_data_0;

  OR2X2 C7788 ( .A(N163), .B(N164), .Y(N165) );
  INVX2 I_25 ( .A(N161), .Y(N162) );
  INVX2 I_23 ( .A(N158), .Y(N159) );
  INVX2 I_22 ( .A(address[3]), .Y(N156) );
  INVX2 I_21 ( .A(N154), .Y(N155) );
  INVX2 I_20 ( .A(N151), .Y(N152) );
  INVX2 I_19 ( .A(address[1]), .Y(N147) );
  INVX2 I_17 ( .A(address[4]), .Y(N141) );
  INVX2 I_16 ( .A(address[5]), .Y(N140) );
  INVX2 I_15 ( .A(address[6]), .Y(N139) );
  INVX2 I_14 ( .A(address[7]), .Y(N138) );
  OR2X2 C7770 ( .A(address[7]), .B(address[6]), .Y(N245) );
  OR2X2 C7769 ( .A(N245), .B(address[5]), .Y(N246) );
  OR2X2 C7768 ( .A(N246), .B(address[4]), .Y(N247) );
  AND2X1 C7767 ( .A(N247), .B(N128), .Y(N129) );
  AND2X1 C7697 ( .A(N199), .B(N212), .Y(N244) );
  AND2X1 C7696 ( .A(N199), .B(N211), .Y(N243) );
  AND2X1 C7695 ( .A(N199), .B(N210), .Y(N242) );
  AND2X1 C7694 ( .A(N199), .B(N209), .Y(N241) );
  AND2X1 C7693 ( .A(N199), .B(N208), .Y(N240) );
  AND2X1 C7692 ( .A(N199), .B(N207), .Y(N239) );
  AND2X1 C7691 ( .A(N199), .B(N206), .Y(N238) );
  AND2X1 C7690 ( .A(N199), .B(N205), .Y(N237) );
  AND2X1 C7689 ( .A(N198), .B(N212), .Y(N236) );
  AND2X1 C7688 ( .A(N198), .B(N211), .Y(N235) );
  AND2X1 C7687 ( .A(N198), .B(N210), .Y(N234) );
  AND2X1 C7686 ( .A(N198), .B(N209), .Y(N233) );
  AND2X1 C7685 ( .A(N198), .B(N208), .Y(N232) );
  AND2X1 C7684 ( .A(N198), .B(N207), .Y(N231) );
  AND2X1 C7683 ( .A(N198), .B(N206), .Y(N230) );
  AND2X1 C7682 ( .A(N198), .B(N205), .Y(N229) );
  AND2X1 C7681 ( .A(N197), .B(N212), .Y(N228) );
  AND2X1 C7680 ( .A(N197), .B(N211), .Y(N227) );
  AND2X1 C7679 ( .A(N197), .B(N210), .Y(N226) );
  AND2X1 C7678 ( .A(N197), .B(N209), .Y(N225) );
  AND2X1 C7677 ( .A(N197), .B(N208), .Y(N224) );
  AND2X1 C7676 ( .A(N197), .B(N207), .Y(N223) );
  AND2X1 C7675 ( .A(N197), .B(N206), .Y(N222) );
  AND2X1 C7674 ( .A(N197), .B(N205), .Y(N221) );
  AND2X1 C7673 ( .A(N196), .B(N212), .Y(N220) );
  AND2X1 C7672 ( .A(N196), .B(N211), .Y(N219) );
  AND2X1 C7671 ( .A(N196), .B(N210), .Y(N218) );
  AND2X1 C7670 ( .A(N196), .B(N209), .Y(N217) );
  AND2X1 C7669 ( .A(N196), .B(N208), .Y(N216) );
  AND2X1 C7668 ( .A(N196), .B(N207), .Y(N215) );
  AND2X1 C7667 ( .A(N196), .B(N206), .Y(N214) );
  AND2X1 C7666 ( .A(N196), .B(N205), .Y(N213) );
  AND2X1 C7665 ( .A(N200), .B(N204), .Y(N212) );
  AND2X1 C7664 ( .A(N200), .B(N203), .Y(N211) );
  AND2X1 C7663 ( .A(N200), .B(N202), .Y(N210) );
  AND2X1 C7662 ( .A(N200), .B(N201), .Y(N209) );
  AND2X1 C7661 ( .A(address[2]), .B(N204), .Y(N208) );
  AND2X1 C7660 ( .A(address[2]), .B(N203), .Y(N207) );
  AND2X1 C7659 ( .A(address[2]), .B(N202), .Y(N206) );
  AND2X1 C7658 ( .A(address[2]), .B(N201), .Y(N205) );
  INVX2 I_8 ( .A(address[1]), .Y(N7) );
  INVX2 I_7 ( .A(address[0]), .Y(N6) );
  AND2X1 C7657 ( .A(N6), .B(N7), .Y(N204) );
  INVX2 I_6 ( .A(address[1]), .Y(N5) );
  AND2X1 C7656 ( .A(address[0]), .B(N5), .Y(N203) );
  INVX2 I_5 ( .A(address[0]), .Y(N4) );
  AND2X1 C7655 ( .A(N4), .B(address[1]), .Y(N202) );
  AND2X1 C7654 ( .A(address[0]), .B(address[1]), .Y(N201) );
  INVX2 I_4 ( .A(address[2]), .Y(N200) );
  INVX2 I_3 ( .A(address[4]), .Y(N3) );
  INVX2 I_2 ( .A(address[3]), .Y(N2) );
  AND2X1 C7652 ( .A(N2), .B(N3), .Y(N199) );
  INVX2 I_1 ( .A(address[4]), .Y(N1) );
  AND2X1 C7651 ( .A(address[3]), .B(N1), .Y(N198) );
  INVX2 I_0 ( .A(address[3]), .Y(N0) );
  AND2X1 C7650 ( .A(N0), .B(address[4]), .Y(N197) );
  AND2X1 C7649 ( .A(address[3]), .B(address[4]), .Y(N196) );
  OR2X2 C7399 ( .A(N156), .B(address[1]), .Y(N157) );
  OR2X2 C7395 ( .A(address[3]), .B(N147), .Y(N153) );
  OR2X2 C7391 ( .A(address[3]), .B(address[1]), .Y(N150) );
  AND2X1 C7388 ( .A(N156), .B(N147), .Y(N148) );
  AND2X1 C7380 ( .A(N142), .B(N143), .Y(N144) );
  AND2X1 C7379 ( .A(N140), .B(N141), .Y(N143) );
  AND2X1 C7378 ( .A(N138), .B(N139), .Y(N142) );
  DFFPOSX1 next_reg_reg ( .D(n2172), .CLK(clk), .Q(core_next) );
  DFFPOSX1 \block_mem_reg[0][31]  ( .D(n2106), .CLK(clk), .Q(core_block[1023])
         );
  DFFPOSX1 \block_mem_reg[0][30]  ( .D(n2105), .CLK(clk), .Q(core_block[1022])
         );
  DFFPOSX1 \block_mem_reg[0][29]  ( .D(n2104), .CLK(clk), .Q(core_block[1021])
         );
  DFFPOSX1 \block_mem_reg[0][28]  ( .D(n2103), .CLK(clk), .Q(core_block[1020])
         );
  DFFPOSX1 \block_mem_reg[0][27]  ( .D(n2102), .CLK(clk), .Q(core_block[1019])
         );
  DFFPOSX1 \block_mem_reg[0][26]  ( .D(n2101), .CLK(clk), .Q(core_block[1018])
         );
  DFFPOSX1 \block_mem_reg[0][25]  ( .D(n2100), .CLK(clk), .Q(core_block[1017])
         );
  DFFPOSX1 \block_mem_reg[0][24]  ( .D(n2099), .CLK(clk), .Q(core_block[1016])
         );
  DFFPOSX1 \block_mem_reg[0][23]  ( .D(n2098), .CLK(clk), .Q(core_block[1015])
         );
  DFFPOSX1 \block_mem_reg[0][22]  ( .D(n2097), .CLK(clk), .Q(core_block[1014])
         );
  DFFPOSX1 \block_mem_reg[0][21]  ( .D(n2096), .CLK(clk), .Q(core_block[1013])
         );
  DFFPOSX1 \block_mem_reg[0][20]  ( .D(n2095), .CLK(clk), .Q(core_block[1012])
         );
  DFFPOSX1 \block_mem_reg[0][19]  ( .D(n2094), .CLK(clk), .Q(core_block[1011])
         );
  DFFPOSX1 \block_mem_reg[0][18]  ( .D(n2093), .CLK(clk), .Q(core_block[1010])
         );
  DFFPOSX1 \block_mem_reg[0][17]  ( .D(n2092), .CLK(clk), .Q(core_block[1009])
         );
  DFFPOSX1 \block_mem_reg[0][16]  ( .D(n2091), .CLK(clk), .Q(core_block[1008])
         );
  DFFPOSX1 \block_mem_reg[0][15]  ( .D(n2090), .CLK(clk), .Q(core_block[1007])
         );
  DFFPOSX1 \block_mem_reg[0][14]  ( .D(n2089), .CLK(clk), .Q(core_block[1006])
         );
  DFFPOSX1 \block_mem_reg[0][13]  ( .D(n2088), .CLK(clk), .Q(core_block[1005])
         );
  DFFPOSX1 \block_mem_reg[0][12]  ( .D(n2087), .CLK(clk), .Q(core_block[1004])
         );
  DFFPOSX1 \block_mem_reg[0][11]  ( .D(n2086), .CLK(clk), .Q(core_block[1003])
         );
  DFFPOSX1 \block_mem_reg[0][10]  ( .D(n2085), .CLK(clk), .Q(core_block[1002])
         );
  DFFPOSX1 \block_mem_reg[0][9]  ( .D(n2084), .CLK(clk), .Q(core_block[1001])
         );
  DFFPOSX1 \block_mem_reg[0][8]  ( .D(n2083), .CLK(clk), .Q(core_block[1000])
         );
  DFFPOSX1 \block_mem_reg[0][7]  ( .D(n2082), .CLK(clk), .Q(core_block[999])
         );
  DFFPOSX1 \block_mem_reg[0][6]  ( .D(n2081), .CLK(clk), .Q(core_block[998])
         );
  DFFPOSX1 \block_mem_reg[0][5]  ( .D(n2080), .CLK(clk), .Q(core_block[997])
         );
  DFFPOSX1 \block_mem_reg[0][4]  ( .D(n2079), .CLK(clk), .Q(core_block[996])
         );
  DFFPOSX1 \block_mem_reg[0][3]  ( .D(n2078), .CLK(clk), .Q(core_block[995])
         );
  DFFPOSX1 \block_mem_reg[0][2]  ( .D(n2077), .CLK(clk), .Q(core_block[994])
         );
  DFFPOSX1 \block_mem_reg[0][1]  ( .D(n2076), .CLK(clk), .Q(core_block[993])
         );
  DFFPOSX1 \block_mem_reg[0][0]  ( .D(n2075), .CLK(clk), .Q(core_block[992])
         );
  DFFPOSX1 \block_mem_reg[1][31]  ( .D(n2074), .CLK(clk), .Q(core_block[991])
         );
  DFFPOSX1 \block_mem_reg[1][30]  ( .D(n2073), .CLK(clk), .Q(core_block[990])
         );
  DFFPOSX1 \block_mem_reg[1][29]  ( .D(n2072), .CLK(clk), .Q(core_block[989])
         );
  DFFPOSX1 \block_mem_reg[1][28]  ( .D(n2071), .CLK(clk), .Q(core_block[988])
         );
  DFFPOSX1 \block_mem_reg[1][27]  ( .D(n2070), .CLK(clk), .Q(core_block[987])
         );
  DFFPOSX1 \block_mem_reg[1][26]  ( .D(n2069), .CLK(clk), .Q(core_block[986])
         );
  DFFPOSX1 \block_mem_reg[1][25]  ( .D(n2068), .CLK(clk), .Q(core_block[985])
         );
  DFFPOSX1 \block_mem_reg[1][24]  ( .D(n2067), .CLK(clk), .Q(core_block[984])
         );
  DFFPOSX1 \block_mem_reg[1][23]  ( .D(n2066), .CLK(clk), .Q(core_block[983])
         );
  DFFPOSX1 \block_mem_reg[1][22]  ( .D(n2065), .CLK(clk), .Q(core_block[982])
         );
  DFFPOSX1 \block_mem_reg[1][21]  ( .D(n2064), .CLK(clk), .Q(core_block[981])
         );
  DFFPOSX1 \block_mem_reg[1][20]  ( .D(n2063), .CLK(clk), .Q(core_block[980])
         );
  DFFPOSX1 \block_mem_reg[1][19]  ( .D(n2062), .CLK(clk), .Q(core_block[979])
         );
  DFFPOSX1 \block_mem_reg[1][18]  ( .D(n2061), .CLK(clk), .Q(core_block[978])
         );
  DFFPOSX1 \block_mem_reg[1][17]  ( .D(n2060), .CLK(clk), .Q(core_block[977])
         );
  DFFPOSX1 \block_mem_reg[1][16]  ( .D(n2059), .CLK(clk), .Q(core_block[976])
         );
  DFFPOSX1 \block_mem_reg[1][15]  ( .D(n2058), .CLK(clk), .Q(core_block[975])
         );
  DFFPOSX1 \block_mem_reg[1][14]  ( .D(n2057), .CLK(clk), .Q(core_block[974])
         );
  DFFPOSX1 \block_mem_reg[1][13]  ( .D(n2056), .CLK(clk), .Q(core_block[973])
         );
  DFFPOSX1 \block_mem_reg[1][12]  ( .D(n2055), .CLK(clk), .Q(core_block[972])
         );
  DFFPOSX1 \block_mem_reg[1][11]  ( .D(n2054), .CLK(clk), .Q(core_block[971])
         );
  DFFPOSX1 \block_mem_reg[1][10]  ( .D(n2053), .CLK(clk), .Q(core_block[970])
         );
  DFFPOSX1 \block_mem_reg[1][9]  ( .D(n2052), .CLK(clk), .Q(core_block[969])
         );
  DFFPOSX1 \block_mem_reg[1][8]  ( .D(n2051), .CLK(clk), .Q(core_block[968])
         );
  DFFPOSX1 \block_mem_reg[1][7]  ( .D(n2050), .CLK(clk), .Q(core_block[967])
         );
  DFFPOSX1 \block_mem_reg[1][6]  ( .D(n2049), .CLK(clk), .Q(core_block[966])
         );
  DFFPOSX1 \block_mem_reg[1][5]  ( .D(n2048), .CLK(clk), .Q(core_block[965])
         );
  DFFPOSX1 \block_mem_reg[1][4]  ( .D(n2047), .CLK(clk), .Q(core_block[964])
         );
  DFFPOSX1 \block_mem_reg[1][3]  ( .D(n2046), .CLK(clk), .Q(core_block[963])
         );
  DFFPOSX1 \block_mem_reg[1][2]  ( .D(n2045), .CLK(clk), .Q(core_block[962])
         );
  DFFPOSX1 \block_mem_reg[1][1]  ( .D(n2044), .CLK(clk), .Q(core_block[961])
         );
  DFFPOSX1 \block_mem_reg[1][0]  ( .D(n2043), .CLK(clk), .Q(core_block[960])
         );
  DFFPOSX1 \block_mem_reg[2][31]  ( .D(n2042), .CLK(clk), .Q(core_block[959])
         );
  DFFPOSX1 \block_mem_reg[2][30]  ( .D(n2041), .CLK(clk), .Q(core_block[958])
         );
  DFFPOSX1 \block_mem_reg[2][29]  ( .D(n2040), .CLK(clk), .Q(core_block[957])
         );
  DFFPOSX1 \block_mem_reg[2][28]  ( .D(n2039), .CLK(clk), .Q(core_block[956])
         );
  DFFPOSX1 \block_mem_reg[2][27]  ( .D(n2038), .CLK(clk), .Q(core_block[955])
         );
  DFFPOSX1 \block_mem_reg[2][26]  ( .D(n2037), .CLK(clk), .Q(core_block[954])
         );
  DFFPOSX1 \block_mem_reg[2][25]  ( .D(n2036), .CLK(clk), .Q(core_block[953])
         );
  DFFPOSX1 \block_mem_reg[2][24]  ( .D(n2035), .CLK(clk), .Q(core_block[952])
         );
  DFFPOSX1 \block_mem_reg[2][23]  ( .D(n2034), .CLK(clk), .Q(core_block[951])
         );
  DFFPOSX1 \block_mem_reg[2][22]  ( .D(n2033), .CLK(clk), .Q(core_block[950])
         );
  DFFPOSX1 \block_mem_reg[2][21]  ( .D(n2032), .CLK(clk), .Q(core_block[949])
         );
  DFFPOSX1 \block_mem_reg[2][20]  ( .D(n2031), .CLK(clk), .Q(core_block[948])
         );
  DFFPOSX1 \block_mem_reg[2][19]  ( .D(n2030), .CLK(clk), .Q(core_block[947])
         );
  DFFPOSX1 \block_mem_reg[2][18]  ( .D(n2029), .CLK(clk), .Q(core_block[946])
         );
  DFFPOSX1 \block_mem_reg[2][17]  ( .D(n2028), .CLK(clk), .Q(core_block[945])
         );
  DFFPOSX1 \block_mem_reg[2][16]  ( .D(n2027), .CLK(clk), .Q(core_block[944])
         );
  DFFPOSX1 \block_mem_reg[2][15]  ( .D(n2026), .CLK(clk), .Q(core_block[943])
         );
  DFFPOSX1 \block_mem_reg[2][14]  ( .D(n2025), .CLK(clk), .Q(core_block[942])
         );
  DFFPOSX1 \block_mem_reg[2][13]  ( .D(n2024), .CLK(clk), .Q(core_block[941])
         );
  DFFPOSX1 \block_mem_reg[2][12]  ( .D(n2023), .CLK(clk), .Q(core_block[940])
         );
  DFFPOSX1 \block_mem_reg[2][11]  ( .D(n2022), .CLK(clk), .Q(core_block[939])
         );
  DFFPOSX1 \block_mem_reg[2][10]  ( .D(n2021), .CLK(clk), .Q(core_block[938])
         );
  DFFPOSX1 \block_mem_reg[2][9]  ( .D(n2020), .CLK(clk), .Q(core_block[937])
         );
  DFFPOSX1 \block_mem_reg[2][8]  ( .D(n2019), .CLK(clk), .Q(core_block[936])
         );
  DFFPOSX1 \block_mem_reg[2][7]  ( .D(n2018), .CLK(clk), .Q(core_block[935])
         );
  DFFPOSX1 \block_mem_reg[2][6]  ( .D(n2017), .CLK(clk), .Q(core_block[934])
         );
  DFFPOSX1 \block_mem_reg[2][5]  ( .D(n2016), .CLK(clk), .Q(core_block[933])
         );
  DFFPOSX1 \block_mem_reg[2][4]  ( .D(n2015), .CLK(clk), .Q(core_block[932])
         );
  DFFPOSX1 \block_mem_reg[2][3]  ( .D(n2014), .CLK(clk), .Q(core_block[931])
         );
  DFFPOSX1 \block_mem_reg[2][2]  ( .D(n2013), .CLK(clk), .Q(core_block[930])
         );
  DFFPOSX1 \block_mem_reg[2][1]  ( .D(n2012), .CLK(clk), .Q(core_block[929])
         );
  DFFPOSX1 \block_mem_reg[2][0]  ( .D(n2011), .CLK(clk), .Q(core_block[928])
         );
  DFFPOSX1 \block_mem_reg[3][31]  ( .D(n2010), .CLK(clk), .Q(core_block[927])
         );
  DFFPOSX1 \block_mem_reg[3][30]  ( .D(n2009), .CLK(clk), .Q(core_block[926])
         );
  DFFPOSX1 \block_mem_reg[3][29]  ( .D(n2008), .CLK(clk), .Q(core_block[925])
         );
  DFFPOSX1 \block_mem_reg[3][28]  ( .D(n2007), .CLK(clk), .Q(core_block[924])
         );
  DFFPOSX1 \block_mem_reg[3][27]  ( .D(n2006), .CLK(clk), .Q(core_block[923])
         );
  DFFPOSX1 \block_mem_reg[3][26]  ( .D(n2005), .CLK(clk), .Q(core_block[922])
         );
  DFFPOSX1 \block_mem_reg[3][25]  ( .D(n2004), .CLK(clk), .Q(core_block[921])
         );
  DFFPOSX1 \block_mem_reg[3][24]  ( .D(n2003), .CLK(clk), .Q(core_block[920])
         );
  DFFPOSX1 \block_mem_reg[3][23]  ( .D(n2002), .CLK(clk), .Q(core_block[919])
         );
  DFFPOSX1 \block_mem_reg[3][22]  ( .D(n2001), .CLK(clk), .Q(core_block[918])
         );
  DFFPOSX1 \block_mem_reg[3][21]  ( .D(n2000), .CLK(clk), .Q(core_block[917])
         );
  DFFPOSX1 \block_mem_reg[3][20]  ( .D(n1999), .CLK(clk), .Q(core_block[916])
         );
  DFFPOSX1 \block_mem_reg[3][19]  ( .D(n1998), .CLK(clk), .Q(core_block[915])
         );
  DFFPOSX1 \block_mem_reg[3][18]  ( .D(n1997), .CLK(clk), .Q(core_block[914])
         );
  DFFPOSX1 \block_mem_reg[3][17]  ( .D(n1996), .CLK(clk), .Q(core_block[913])
         );
  DFFPOSX1 \block_mem_reg[3][16]  ( .D(n1995), .CLK(clk), .Q(core_block[912])
         );
  DFFPOSX1 \block_mem_reg[3][15]  ( .D(n1994), .CLK(clk), .Q(core_block[911])
         );
  DFFPOSX1 \block_mem_reg[3][14]  ( .D(n1993), .CLK(clk), .Q(core_block[910])
         );
  DFFPOSX1 \block_mem_reg[3][13]  ( .D(n1992), .CLK(clk), .Q(core_block[909])
         );
  DFFPOSX1 \block_mem_reg[3][12]  ( .D(n1991), .CLK(clk), .Q(core_block[908])
         );
  DFFPOSX1 \block_mem_reg[3][11]  ( .D(n1990), .CLK(clk), .Q(core_block[907])
         );
  DFFPOSX1 \block_mem_reg[3][10]  ( .D(n1989), .CLK(clk), .Q(core_block[906])
         );
  DFFPOSX1 \block_mem_reg[3][9]  ( .D(n1988), .CLK(clk), .Q(core_block[905])
         );
  DFFPOSX1 \block_mem_reg[3][8]  ( .D(n1987), .CLK(clk), .Q(core_block[904])
         );
  DFFPOSX1 \block_mem_reg[3][7]  ( .D(n1986), .CLK(clk), .Q(core_block[903])
         );
  DFFPOSX1 \block_mem_reg[3][6]  ( .D(n1985), .CLK(clk), .Q(core_block[902])
         );
  DFFPOSX1 \block_mem_reg[3][5]  ( .D(n1984), .CLK(clk), .Q(core_block[901])
         );
  DFFPOSX1 \block_mem_reg[3][4]  ( .D(n1983), .CLK(clk), .Q(core_block[900])
         );
  DFFPOSX1 \block_mem_reg[3][3]  ( .D(n1982), .CLK(clk), .Q(core_block[899])
         );
  DFFPOSX1 \block_mem_reg[3][2]  ( .D(n1981), .CLK(clk), .Q(core_block[898])
         );
  DFFPOSX1 \block_mem_reg[3][1]  ( .D(n1980), .CLK(clk), .Q(core_block[897])
         );
  DFFPOSX1 \block_mem_reg[3][0]  ( .D(n1979), .CLK(clk), .Q(core_block[896])
         );
  DFFPOSX1 \block_mem_reg[4][31]  ( .D(n1978), .CLK(clk), .Q(core_block[895])
         );
  DFFPOSX1 \block_mem_reg[4][30]  ( .D(n1977), .CLK(clk), .Q(core_block[894])
         );
  DFFPOSX1 \block_mem_reg[4][29]  ( .D(n1976), .CLK(clk), .Q(core_block[893])
         );
  DFFPOSX1 \block_mem_reg[4][28]  ( .D(n1975), .CLK(clk), .Q(core_block[892])
         );
  DFFPOSX1 \block_mem_reg[4][27]  ( .D(n1974), .CLK(clk), .Q(core_block[891])
         );
  DFFPOSX1 \block_mem_reg[4][26]  ( .D(n1973), .CLK(clk), .Q(core_block[890])
         );
  DFFPOSX1 \block_mem_reg[4][25]  ( .D(n1972), .CLK(clk), .Q(core_block[889])
         );
  DFFPOSX1 \block_mem_reg[4][24]  ( .D(n1971), .CLK(clk), .Q(core_block[888])
         );
  DFFPOSX1 \block_mem_reg[4][23]  ( .D(n1970), .CLK(clk), .Q(core_block[887])
         );
  DFFPOSX1 \block_mem_reg[4][22]  ( .D(n1969), .CLK(clk), .Q(core_block[886])
         );
  DFFPOSX1 \block_mem_reg[4][21]  ( .D(n1968), .CLK(clk), .Q(core_block[885])
         );
  DFFPOSX1 \block_mem_reg[4][20]  ( .D(n1967), .CLK(clk), .Q(core_block[884])
         );
  DFFPOSX1 \block_mem_reg[4][19]  ( .D(n1966), .CLK(clk), .Q(core_block[883])
         );
  DFFPOSX1 \block_mem_reg[4][18]  ( .D(n1965), .CLK(clk), .Q(core_block[882])
         );
  DFFPOSX1 \block_mem_reg[4][17]  ( .D(n1964), .CLK(clk), .Q(core_block[881])
         );
  DFFPOSX1 \block_mem_reg[4][16]  ( .D(n1963), .CLK(clk), .Q(core_block[880])
         );
  DFFPOSX1 \block_mem_reg[4][15]  ( .D(n1962), .CLK(clk), .Q(core_block[879])
         );
  DFFPOSX1 \block_mem_reg[4][14]  ( .D(n1961), .CLK(clk), .Q(core_block[878])
         );
  DFFPOSX1 \block_mem_reg[4][13]  ( .D(n1960), .CLK(clk), .Q(core_block[877])
         );
  DFFPOSX1 \block_mem_reg[4][12]  ( .D(n1959), .CLK(clk), .Q(core_block[876])
         );
  DFFPOSX1 \block_mem_reg[4][11]  ( .D(n1958), .CLK(clk), .Q(core_block[875])
         );
  DFFPOSX1 \block_mem_reg[4][10]  ( .D(n1957), .CLK(clk), .Q(core_block[874])
         );
  DFFPOSX1 \block_mem_reg[4][9]  ( .D(n1956), .CLK(clk), .Q(core_block[873])
         );
  DFFPOSX1 \block_mem_reg[4][8]  ( .D(n1955), .CLK(clk), .Q(core_block[872])
         );
  DFFPOSX1 \block_mem_reg[4][7]  ( .D(n1954), .CLK(clk), .Q(core_block[871])
         );
  DFFPOSX1 \block_mem_reg[4][6]  ( .D(n1953), .CLK(clk), .Q(core_block[870])
         );
  DFFPOSX1 \block_mem_reg[4][5]  ( .D(n1952), .CLK(clk), .Q(core_block[869])
         );
  DFFPOSX1 \block_mem_reg[4][4]  ( .D(n1951), .CLK(clk), .Q(core_block[868])
         );
  DFFPOSX1 \block_mem_reg[4][3]  ( .D(n1950), .CLK(clk), .Q(core_block[867])
         );
  DFFPOSX1 \block_mem_reg[4][2]  ( .D(n1949), .CLK(clk), .Q(core_block[866])
         );
  DFFPOSX1 \block_mem_reg[4][1]  ( .D(n1948), .CLK(clk), .Q(core_block[865])
         );
  DFFPOSX1 \block_mem_reg[4][0]  ( .D(n1947), .CLK(clk), .Q(core_block[864])
         );
  DFFPOSX1 \block_mem_reg[5][31]  ( .D(n1946), .CLK(clk), .Q(core_block[863])
         );
  DFFPOSX1 \block_mem_reg[5][30]  ( .D(n1945), .CLK(clk), .Q(core_block[862])
         );
  DFFPOSX1 \block_mem_reg[5][29]  ( .D(n1944), .CLK(clk), .Q(core_block[861])
         );
  DFFPOSX1 \block_mem_reg[5][28]  ( .D(n1943), .CLK(clk), .Q(core_block[860])
         );
  DFFPOSX1 \block_mem_reg[5][27]  ( .D(n1942), .CLK(clk), .Q(core_block[859])
         );
  DFFPOSX1 \block_mem_reg[5][26]  ( .D(n1941), .CLK(clk), .Q(core_block[858])
         );
  DFFPOSX1 \block_mem_reg[5][25]  ( .D(n1940), .CLK(clk), .Q(core_block[857])
         );
  DFFPOSX1 \block_mem_reg[5][24]  ( .D(n1939), .CLK(clk), .Q(core_block[856])
         );
  DFFPOSX1 \block_mem_reg[5][23]  ( .D(n1938), .CLK(clk), .Q(core_block[855])
         );
  DFFPOSX1 \block_mem_reg[5][22]  ( .D(n1937), .CLK(clk), .Q(core_block[854])
         );
  DFFPOSX1 \block_mem_reg[5][21]  ( .D(n1936), .CLK(clk), .Q(core_block[853])
         );
  DFFPOSX1 \block_mem_reg[5][20]  ( .D(n1935), .CLK(clk), .Q(core_block[852])
         );
  DFFPOSX1 \block_mem_reg[5][19]  ( .D(n1934), .CLK(clk), .Q(core_block[851])
         );
  DFFPOSX1 \block_mem_reg[5][18]  ( .D(n1933), .CLK(clk), .Q(core_block[850])
         );
  DFFPOSX1 \block_mem_reg[5][17]  ( .D(n1932), .CLK(clk), .Q(core_block[849])
         );
  DFFPOSX1 \block_mem_reg[5][16]  ( .D(n1931), .CLK(clk), .Q(core_block[848])
         );
  DFFPOSX1 \block_mem_reg[5][15]  ( .D(n1930), .CLK(clk), .Q(core_block[847])
         );
  DFFPOSX1 \block_mem_reg[5][14]  ( .D(n1929), .CLK(clk), .Q(core_block[846])
         );
  DFFPOSX1 \block_mem_reg[5][13]  ( .D(n1928), .CLK(clk), .Q(core_block[845])
         );
  DFFPOSX1 \block_mem_reg[5][12]  ( .D(n1927), .CLK(clk), .Q(core_block[844])
         );
  DFFPOSX1 \block_mem_reg[5][11]  ( .D(n1926), .CLK(clk), .Q(core_block[843])
         );
  DFFPOSX1 \block_mem_reg[5][10]  ( .D(n1925), .CLK(clk), .Q(core_block[842])
         );
  DFFPOSX1 \block_mem_reg[5][9]  ( .D(n1924), .CLK(clk), .Q(core_block[841])
         );
  DFFPOSX1 \block_mem_reg[5][8]  ( .D(n1923), .CLK(clk), .Q(core_block[840])
         );
  DFFPOSX1 \block_mem_reg[5][7]  ( .D(n1922), .CLK(clk), .Q(core_block[839])
         );
  DFFPOSX1 \block_mem_reg[5][6]  ( .D(n1921), .CLK(clk), .Q(core_block[838])
         );
  DFFPOSX1 \block_mem_reg[5][5]  ( .D(n1920), .CLK(clk), .Q(core_block[837])
         );
  DFFPOSX1 \block_mem_reg[5][4]  ( .D(n1919), .CLK(clk), .Q(core_block[836])
         );
  DFFPOSX1 \block_mem_reg[5][3]  ( .D(n1918), .CLK(clk), .Q(core_block[835])
         );
  DFFPOSX1 \block_mem_reg[5][2]  ( .D(n1917), .CLK(clk), .Q(core_block[834])
         );
  DFFPOSX1 \block_mem_reg[5][1]  ( .D(n1916), .CLK(clk), .Q(core_block[833])
         );
  DFFPOSX1 \block_mem_reg[5][0]  ( .D(n1915), .CLK(clk), .Q(core_block[832])
         );
  DFFPOSX1 \block_mem_reg[6][31]  ( .D(n1914), .CLK(clk), .Q(core_block[831])
         );
  DFFPOSX1 \block_mem_reg[6][30]  ( .D(n1913), .CLK(clk), .Q(core_block[830])
         );
  DFFPOSX1 \block_mem_reg[6][29]  ( .D(n1912), .CLK(clk), .Q(core_block[829])
         );
  DFFPOSX1 \block_mem_reg[6][28]  ( .D(n1911), .CLK(clk), .Q(core_block[828])
         );
  DFFPOSX1 \block_mem_reg[6][27]  ( .D(n1910), .CLK(clk), .Q(core_block[827])
         );
  DFFPOSX1 \block_mem_reg[6][26]  ( .D(n1909), .CLK(clk), .Q(core_block[826])
         );
  DFFPOSX1 \block_mem_reg[6][25]  ( .D(n1908), .CLK(clk), .Q(core_block[825])
         );
  DFFPOSX1 \block_mem_reg[6][24]  ( .D(n1907), .CLK(clk), .Q(core_block[824])
         );
  DFFPOSX1 \block_mem_reg[6][23]  ( .D(n1906), .CLK(clk), .Q(core_block[823])
         );
  DFFPOSX1 \block_mem_reg[6][22]  ( .D(n1905), .CLK(clk), .Q(core_block[822])
         );
  DFFPOSX1 \block_mem_reg[6][21]  ( .D(n1904), .CLK(clk), .Q(core_block[821])
         );
  DFFPOSX1 \block_mem_reg[6][20]  ( .D(n1903), .CLK(clk), .Q(core_block[820])
         );
  DFFPOSX1 \block_mem_reg[6][19]  ( .D(n1902), .CLK(clk), .Q(core_block[819])
         );
  DFFPOSX1 \block_mem_reg[6][18]  ( .D(n1901), .CLK(clk), .Q(core_block[818])
         );
  DFFPOSX1 \block_mem_reg[6][17]  ( .D(n1900), .CLK(clk), .Q(core_block[817])
         );
  DFFPOSX1 \block_mem_reg[6][16]  ( .D(n1899), .CLK(clk), .Q(core_block[816])
         );
  DFFPOSX1 \block_mem_reg[6][15]  ( .D(n1898), .CLK(clk), .Q(core_block[815])
         );
  DFFPOSX1 \block_mem_reg[6][14]  ( .D(n1897), .CLK(clk), .Q(core_block[814])
         );
  DFFPOSX1 \block_mem_reg[6][13]  ( .D(n1896), .CLK(clk), .Q(core_block[813])
         );
  DFFPOSX1 \block_mem_reg[6][12]  ( .D(n1895), .CLK(clk), .Q(core_block[812])
         );
  DFFPOSX1 \block_mem_reg[6][11]  ( .D(n1894), .CLK(clk), .Q(core_block[811])
         );
  DFFPOSX1 \block_mem_reg[6][10]  ( .D(n1893), .CLK(clk), .Q(core_block[810])
         );
  DFFPOSX1 \block_mem_reg[6][9]  ( .D(n1892), .CLK(clk), .Q(core_block[809])
         );
  DFFPOSX1 \block_mem_reg[6][8]  ( .D(n1891), .CLK(clk), .Q(core_block[808])
         );
  DFFPOSX1 \block_mem_reg[6][7]  ( .D(n1890), .CLK(clk), .Q(core_block[807])
         );
  DFFPOSX1 \block_mem_reg[6][6]  ( .D(n1889), .CLK(clk), .Q(core_block[806])
         );
  DFFPOSX1 \block_mem_reg[6][5]  ( .D(n1888), .CLK(clk), .Q(core_block[805])
         );
  DFFPOSX1 \block_mem_reg[6][4]  ( .D(n1887), .CLK(clk), .Q(core_block[804])
         );
  DFFPOSX1 \block_mem_reg[6][3]  ( .D(n1886), .CLK(clk), .Q(core_block[803])
         );
  DFFPOSX1 \block_mem_reg[6][2]  ( .D(n1885), .CLK(clk), .Q(core_block[802])
         );
  DFFPOSX1 \block_mem_reg[6][1]  ( .D(n1884), .CLK(clk), .Q(core_block[801])
         );
  DFFPOSX1 \block_mem_reg[6][0]  ( .D(n1883), .CLK(clk), .Q(core_block[800])
         );
  DFFPOSX1 \block_mem_reg[7][31]  ( .D(n1882), .CLK(clk), .Q(core_block[799])
         );
  DFFPOSX1 \block_mem_reg[7][30]  ( .D(n1881), .CLK(clk), .Q(core_block[798])
         );
  DFFPOSX1 \block_mem_reg[7][29]  ( .D(n1880), .CLK(clk), .Q(core_block[797])
         );
  DFFPOSX1 \block_mem_reg[7][28]  ( .D(n1879), .CLK(clk), .Q(core_block[796])
         );
  DFFPOSX1 \block_mem_reg[7][27]  ( .D(n1878), .CLK(clk), .Q(core_block[795])
         );
  DFFPOSX1 \block_mem_reg[7][26]  ( .D(n1877), .CLK(clk), .Q(core_block[794])
         );
  DFFPOSX1 \block_mem_reg[7][25]  ( .D(n1876), .CLK(clk), .Q(core_block[793])
         );
  DFFPOSX1 \block_mem_reg[7][24]  ( .D(n1875), .CLK(clk), .Q(core_block[792])
         );
  DFFPOSX1 \block_mem_reg[7][23]  ( .D(n1874), .CLK(clk), .Q(core_block[791])
         );
  DFFPOSX1 \block_mem_reg[7][22]  ( .D(n1873), .CLK(clk), .Q(core_block[790])
         );
  DFFPOSX1 \block_mem_reg[7][21]  ( .D(n1872), .CLK(clk), .Q(core_block[789])
         );
  DFFPOSX1 \block_mem_reg[7][20]  ( .D(n1871), .CLK(clk), .Q(core_block[788])
         );
  DFFPOSX1 \block_mem_reg[7][19]  ( .D(n1870), .CLK(clk), .Q(core_block[787])
         );
  DFFPOSX1 \block_mem_reg[7][18]  ( .D(n1869), .CLK(clk), .Q(core_block[786])
         );
  DFFPOSX1 \block_mem_reg[7][17]  ( .D(n1868), .CLK(clk), .Q(core_block[785])
         );
  DFFPOSX1 \block_mem_reg[7][16]  ( .D(n1867), .CLK(clk), .Q(core_block[784])
         );
  DFFPOSX1 \block_mem_reg[7][15]  ( .D(n1866), .CLK(clk), .Q(core_block[783])
         );
  DFFPOSX1 \block_mem_reg[7][14]  ( .D(n1865), .CLK(clk), .Q(core_block[782])
         );
  DFFPOSX1 \block_mem_reg[7][13]  ( .D(n1864), .CLK(clk), .Q(core_block[781])
         );
  DFFPOSX1 \block_mem_reg[7][12]  ( .D(n1863), .CLK(clk), .Q(core_block[780])
         );
  DFFPOSX1 \block_mem_reg[7][11]  ( .D(n1862), .CLK(clk), .Q(core_block[779])
         );
  DFFPOSX1 \block_mem_reg[7][10]  ( .D(n1861), .CLK(clk), .Q(core_block[778])
         );
  DFFPOSX1 \block_mem_reg[7][9]  ( .D(n1860), .CLK(clk), .Q(core_block[777])
         );
  DFFPOSX1 \block_mem_reg[7][8]  ( .D(n1859), .CLK(clk), .Q(core_block[776])
         );
  DFFPOSX1 \block_mem_reg[7][7]  ( .D(n1858), .CLK(clk), .Q(core_block[775])
         );
  DFFPOSX1 \block_mem_reg[7][6]  ( .D(n1857), .CLK(clk), .Q(core_block[774])
         );
  DFFPOSX1 \block_mem_reg[7][5]  ( .D(n1856), .CLK(clk), .Q(core_block[773])
         );
  DFFPOSX1 \block_mem_reg[7][4]  ( .D(n1855), .CLK(clk), .Q(core_block[772])
         );
  DFFPOSX1 \block_mem_reg[7][3]  ( .D(n1854), .CLK(clk), .Q(core_block[771])
         );
  DFFPOSX1 \block_mem_reg[7][2]  ( .D(n1853), .CLK(clk), .Q(core_block[770])
         );
  DFFPOSX1 \block_mem_reg[7][1]  ( .D(n1852), .CLK(clk), .Q(core_block[769])
         );
  DFFPOSX1 \block_mem_reg[7][0]  ( .D(n1851), .CLK(clk), .Q(core_block[768])
         );
  DFFPOSX1 \block_mem_reg[8][31]  ( .D(n1850), .CLK(clk), .Q(core_block[767])
         );
  DFFPOSX1 \block_mem_reg[8][30]  ( .D(n1849), .CLK(clk), .Q(core_block[766])
         );
  DFFPOSX1 \block_mem_reg[8][29]  ( .D(n1848), .CLK(clk), .Q(core_block[765])
         );
  DFFPOSX1 \block_mem_reg[8][28]  ( .D(n1847), .CLK(clk), .Q(core_block[764])
         );
  DFFPOSX1 \block_mem_reg[8][27]  ( .D(n1846), .CLK(clk), .Q(core_block[763])
         );
  DFFPOSX1 \block_mem_reg[8][26]  ( .D(n1845), .CLK(clk), .Q(core_block[762])
         );
  DFFPOSX1 \block_mem_reg[8][25]  ( .D(n1844), .CLK(clk), .Q(core_block[761])
         );
  DFFPOSX1 \block_mem_reg[8][24]  ( .D(n1843), .CLK(clk), .Q(core_block[760])
         );
  DFFPOSX1 \block_mem_reg[8][23]  ( .D(n1842), .CLK(clk), .Q(core_block[759])
         );
  DFFPOSX1 \block_mem_reg[8][22]  ( .D(n1841), .CLK(clk), .Q(core_block[758])
         );
  DFFPOSX1 \block_mem_reg[8][21]  ( .D(n1840), .CLK(clk), .Q(core_block[757])
         );
  DFFPOSX1 \block_mem_reg[8][20]  ( .D(n1839), .CLK(clk), .Q(core_block[756])
         );
  DFFPOSX1 \block_mem_reg[8][19]  ( .D(n1838), .CLK(clk), .Q(core_block[755])
         );
  DFFPOSX1 \block_mem_reg[8][18]  ( .D(n1837), .CLK(clk), .Q(core_block[754])
         );
  DFFPOSX1 \block_mem_reg[8][17]  ( .D(n1836), .CLK(clk), .Q(core_block[753])
         );
  DFFPOSX1 \block_mem_reg[8][16]  ( .D(n1835), .CLK(clk), .Q(core_block[752])
         );
  DFFPOSX1 \block_mem_reg[8][15]  ( .D(n1834), .CLK(clk), .Q(core_block[751])
         );
  DFFPOSX1 \block_mem_reg[8][14]  ( .D(n1833), .CLK(clk), .Q(core_block[750])
         );
  DFFPOSX1 \block_mem_reg[8][13]  ( .D(n1832), .CLK(clk), .Q(core_block[749])
         );
  DFFPOSX1 \block_mem_reg[8][12]  ( .D(n1831), .CLK(clk), .Q(core_block[748])
         );
  DFFPOSX1 \block_mem_reg[8][11]  ( .D(n1830), .CLK(clk), .Q(core_block[747])
         );
  DFFPOSX1 \block_mem_reg[8][10]  ( .D(n1829), .CLK(clk), .Q(core_block[746])
         );
  DFFPOSX1 \block_mem_reg[8][9]  ( .D(n1828), .CLK(clk), .Q(core_block[745])
         );
  DFFPOSX1 \block_mem_reg[8][8]  ( .D(n1827), .CLK(clk), .Q(core_block[744])
         );
  DFFPOSX1 \block_mem_reg[8][7]  ( .D(n1826), .CLK(clk), .Q(core_block[743])
         );
  DFFPOSX1 \block_mem_reg[8][6]  ( .D(n1825), .CLK(clk), .Q(core_block[742])
         );
  DFFPOSX1 \block_mem_reg[8][5]  ( .D(n1824), .CLK(clk), .Q(core_block[741])
         );
  DFFPOSX1 \block_mem_reg[8][4]  ( .D(n1823), .CLK(clk), .Q(core_block[740])
         );
  DFFPOSX1 \block_mem_reg[8][3]  ( .D(n1822), .CLK(clk), .Q(core_block[739])
         );
  DFFPOSX1 \block_mem_reg[8][2]  ( .D(n1821), .CLK(clk), .Q(core_block[738])
         );
  DFFPOSX1 \block_mem_reg[8][1]  ( .D(n1820), .CLK(clk), .Q(core_block[737])
         );
  DFFPOSX1 \block_mem_reg[8][0]  ( .D(n1819), .CLK(clk), .Q(core_block[736])
         );
  DFFPOSX1 \block_mem_reg[9][31]  ( .D(n1818), .CLK(clk), .Q(core_block[735])
         );
  DFFPOSX1 \block_mem_reg[9][30]  ( .D(n1817), .CLK(clk), .Q(core_block[734])
         );
  DFFPOSX1 \block_mem_reg[9][29]  ( .D(n1816), .CLK(clk), .Q(core_block[733])
         );
  DFFPOSX1 \block_mem_reg[9][28]  ( .D(n1815), .CLK(clk), .Q(core_block[732])
         );
  DFFPOSX1 \block_mem_reg[9][27]  ( .D(n1814), .CLK(clk), .Q(core_block[731])
         );
  DFFPOSX1 \block_mem_reg[9][26]  ( .D(n1813), .CLK(clk), .Q(core_block[730])
         );
  DFFPOSX1 \block_mem_reg[9][25]  ( .D(n1812), .CLK(clk), .Q(core_block[729])
         );
  DFFPOSX1 \block_mem_reg[9][24]  ( .D(n1811), .CLK(clk), .Q(core_block[728])
         );
  DFFPOSX1 \block_mem_reg[9][23]  ( .D(n1810), .CLK(clk), .Q(core_block[727])
         );
  DFFPOSX1 \block_mem_reg[9][22]  ( .D(n1809), .CLK(clk), .Q(core_block[726])
         );
  DFFPOSX1 \block_mem_reg[9][21]  ( .D(n1808), .CLK(clk), .Q(core_block[725])
         );
  DFFPOSX1 \block_mem_reg[9][20]  ( .D(n1807), .CLK(clk), .Q(core_block[724])
         );
  DFFPOSX1 \block_mem_reg[9][19]  ( .D(n1806), .CLK(clk), .Q(core_block[723])
         );
  DFFPOSX1 \block_mem_reg[9][18]  ( .D(n1805), .CLK(clk), .Q(core_block[722])
         );
  DFFPOSX1 \block_mem_reg[9][17]  ( .D(n1804), .CLK(clk), .Q(core_block[721])
         );
  DFFPOSX1 \block_mem_reg[9][16]  ( .D(n1803), .CLK(clk), .Q(core_block[720])
         );
  DFFPOSX1 \block_mem_reg[9][15]  ( .D(n1802), .CLK(clk), .Q(core_block[719])
         );
  DFFPOSX1 \block_mem_reg[9][14]  ( .D(n1801), .CLK(clk), .Q(core_block[718])
         );
  DFFPOSX1 \block_mem_reg[9][13]  ( .D(n1800), .CLK(clk), .Q(core_block[717])
         );
  DFFPOSX1 \block_mem_reg[9][12]  ( .D(n1799), .CLK(clk), .Q(core_block[716])
         );
  DFFPOSX1 \block_mem_reg[9][11]  ( .D(n1798), .CLK(clk), .Q(core_block[715])
         );
  DFFPOSX1 \block_mem_reg[9][10]  ( .D(n1797), .CLK(clk), .Q(core_block[714])
         );
  DFFPOSX1 \block_mem_reg[9][9]  ( .D(n1796), .CLK(clk), .Q(core_block[713])
         );
  DFFPOSX1 \block_mem_reg[9][8]  ( .D(n1795), .CLK(clk), .Q(core_block[712])
         );
  DFFPOSX1 \block_mem_reg[9][7]  ( .D(n1794), .CLK(clk), .Q(core_block[711])
         );
  DFFPOSX1 \block_mem_reg[9][6]  ( .D(n1793), .CLK(clk), .Q(core_block[710])
         );
  DFFPOSX1 \block_mem_reg[9][5]  ( .D(n1792), .CLK(clk), .Q(core_block[709])
         );
  DFFPOSX1 \block_mem_reg[9][4]  ( .D(n1791), .CLK(clk), .Q(core_block[708])
         );
  DFFPOSX1 \block_mem_reg[9][3]  ( .D(n1790), .CLK(clk), .Q(core_block[707])
         );
  DFFPOSX1 \block_mem_reg[9][2]  ( .D(n1789), .CLK(clk), .Q(core_block[706])
         );
  DFFPOSX1 \block_mem_reg[9][1]  ( .D(n1788), .CLK(clk), .Q(core_block[705])
         );
  DFFPOSX1 \block_mem_reg[9][0]  ( .D(n1787), .CLK(clk), .Q(core_block[704])
         );
  DFFPOSX1 \block_mem_reg[10][31]  ( .D(n1786), .CLK(clk), .Q(core_block[703])
         );
  DFFPOSX1 \block_mem_reg[10][30]  ( .D(n1785), .CLK(clk), .Q(core_block[702])
         );
  DFFPOSX1 \block_mem_reg[10][29]  ( .D(n1784), .CLK(clk), .Q(core_block[701])
         );
  DFFPOSX1 \block_mem_reg[10][28]  ( .D(n1783), .CLK(clk), .Q(core_block[700])
         );
  DFFPOSX1 \block_mem_reg[10][27]  ( .D(n1782), .CLK(clk), .Q(core_block[699])
         );
  DFFPOSX1 \block_mem_reg[10][26]  ( .D(n1781), .CLK(clk), .Q(core_block[698])
         );
  DFFPOSX1 \block_mem_reg[10][25]  ( .D(n1780), .CLK(clk), .Q(core_block[697])
         );
  DFFPOSX1 \block_mem_reg[10][24]  ( .D(n1779), .CLK(clk), .Q(core_block[696])
         );
  DFFPOSX1 \block_mem_reg[10][23]  ( .D(n1778), .CLK(clk), .Q(core_block[695])
         );
  DFFPOSX1 \block_mem_reg[10][22]  ( .D(n1777), .CLK(clk), .Q(core_block[694])
         );
  DFFPOSX1 \block_mem_reg[10][21]  ( .D(n1776), .CLK(clk), .Q(core_block[693])
         );
  DFFPOSX1 \block_mem_reg[10][20]  ( .D(n1775), .CLK(clk), .Q(core_block[692])
         );
  DFFPOSX1 \block_mem_reg[10][19]  ( .D(n1774), .CLK(clk), .Q(core_block[691])
         );
  DFFPOSX1 \block_mem_reg[10][18]  ( .D(n1773), .CLK(clk), .Q(core_block[690])
         );
  DFFPOSX1 \block_mem_reg[10][17]  ( .D(n1772), .CLK(clk), .Q(core_block[689])
         );
  DFFPOSX1 \block_mem_reg[10][16]  ( .D(n1771), .CLK(clk), .Q(core_block[688])
         );
  DFFPOSX1 \block_mem_reg[10][15]  ( .D(n1770), .CLK(clk), .Q(core_block[687])
         );
  DFFPOSX1 \block_mem_reg[10][14]  ( .D(n1769), .CLK(clk), .Q(core_block[686])
         );
  DFFPOSX1 \block_mem_reg[10][13]  ( .D(n1768), .CLK(clk), .Q(core_block[685])
         );
  DFFPOSX1 \block_mem_reg[10][12]  ( .D(n1767), .CLK(clk), .Q(core_block[684])
         );
  DFFPOSX1 \block_mem_reg[10][11]  ( .D(n1766), .CLK(clk), .Q(core_block[683])
         );
  DFFPOSX1 \block_mem_reg[10][10]  ( .D(n1765), .CLK(clk), .Q(core_block[682])
         );
  DFFPOSX1 \block_mem_reg[10][9]  ( .D(n1764), .CLK(clk), .Q(core_block[681])
         );
  DFFPOSX1 \block_mem_reg[10][8]  ( .D(n1763), .CLK(clk), .Q(core_block[680])
         );
  DFFPOSX1 \block_mem_reg[10][7]  ( .D(n1762), .CLK(clk), .Q(core_block[679])
         );
  DFFPOSX1 \block_mem_reg[10][6]  ( .D(n1761), .CLK(clk), .Q(core_block[678])
         );
  DFFPOSX1 \block_mem_reg[10][5]  ( .D(n1760), .CLK(clk), .Q(core_block[677])
         );
  DFFPOSX1 \block_mem_reg[10][4]  ( .D(n1759), .CLK(clk), .Q(core_block[676])
         );
  DFFPOSX1 \block_mem_reg[10][3]  ( .D(n1758), .CLK(clk), .Q(core_block[675])
         );
  DFFPOSX1 \block_mem_reg[10][2]  ( .D(n1757), .CLK(clk), .Q(core_block[674])
         );
  DFFPOSX1 \block_mem_reg[10][1]  ( .D(n1756), .CLK(clk), .Q(core_block[673])
         );
  DFFPOSX1 \block_mem_reg[10][0]  ( .D(n1755), .CLK(clk), .Q(core_block[672])
         );
  DFFPOSX1 \block_mem_reg[11][31]  ( .D(n1754), .CLK(clk), .Q(core_block[671])
         );
  DFFPOSX1 \block_mem_reg[11][30]  ( .D(n1753), .CLK(clk), .Q(core_block[670])
         );
  DFFPOSX1 \block_mem_reg[11][29]  ( .D(n1752), .CLK(clk), .Q(core_block[669])
         );
  DFFPOSX1 \block_mem_reg[11][28]  ( .D(n1751), .CLK(clk), .Q(core_block[668])
         );
  DFFPOSX1 \block_mem_reg[11][27]  ( .D(n1750), .CLK(clk), .Q(core_block[667])
         );
  DFFPOSX1 \block_mem_reg[11][26]  ( .D(n1749), .CLK(clk), .Q(core_block[666])
         );
  DFFPOSX1 \block_mem_reg[11][25]  ( .D(n1748), .CLK(clk), .Q(core_block[665])
         );
  DFFPOSX1 \block_mem_reg[11][24]  ( .D(n1747), .CLK(clk), .Q(core_block[664])
         );
  DFFPOSX1 \block_mem_reg[11][23]  ( .D(n1746), .CLK(clk), .Q(core_block[663])
         );
  DFFPOSX1 \block_mem_reg[11][22]  ( .D(n1745), .CLK(clk), .Q(core_block[662])
         );
  DFFPOSX1 \block_mem_reg[11][21]  ( .D(n1744), .CLK(clk), .Q(core_block[661])
         );
  DFFPOSX1 \block_mem_reg[11][20]  ( .D(n1743), .CLK(clk), .Q(core_block[660])
         );
  DFFPOSX1 \block_mem_reg[11][19]  ( .D(n1742), .CLK(clk), .Q(core_block[659])
         );
  DFFPOSX1 \block_mem_reg[11][18]  ( .D(n1741), .CLK(clk), .Q(core_block[658])
         );
  DFFPOSX1 \block_mem_reg[11][17]  ( .D(n1740), .CLK(clk), .Q(core_block[657])
         );
  DFFPOSX1 \block_mem_reg[11][16]  ( .D(n1739), .CLK(clk), .Q(core_block[656])
         );
  DFFPOSX1 \block_mem_reg[11][15]  ( .D(n1738), .CLK(clk), .Q(core_block[655])
         );
  DFFPOSX1 \block_mem_reg[11][14]  ( .D(n1737), .CLK(clk), .Q(core_block[654])
         );
  DFFPOSX1 \block_mem_reg[11][13]  ( .D(n1736), .CLK(clk), .Q(core_block[653])
         );
  DFFPOSX1 \block_mem_reg[11][12]  ( .D(n1735), .CLK(clk), .Q(core_block[652])
         );
  DFFPOSX1 \block_mem_reg[11][11]  ( .D(n1734), .CLK(clk), .Q(core_block[651])
         );
  DFFPOSX1 \block_mem_reg[11][10]  ( .D(n1733), .CLK(clk), .Q(core_block[650])
         );
  DFFPOSX1 \block_mem_reg[11][9]  ( .D(n1732), .CLK(clk), .Q(core_block[649])
         );
  DFFPOSX1 \block_mem_reg[11][8]  ( .D(n1731), .CLK(clk), .Q(core_block[648])
         );
  DFFPOSX1 \block_mem_reg[11][7]  ( .D(n1730), .CLK(clk), .Q(core_block[647])
         );
  DFFPOSX1 \block_mem_reg[11][6]  ( .D(n1729), .CLK(clk), .Q(core_block[646])
         );
  DFFPOSX1 \block_mem_reg[11][5]  ( .D(n1728), .CLK(clk), .Q(core_block[645])
         );
  DFFPOSX1 \block_mem_reg[11][4]  ( .D(n1727), .CLK(clk), .Q(core_block[644])
         );
  DFFPOSX1 \block_mem_reg[11][3]  ( .D(n1726), .CLK(clk), .Q(core_block[643])
         );
  DFFPOSX1 \block_mem_reg[11][2]  ( .D(n1725), .CLK(clk), .Q(core_block[642])
         );
  DFFPOSX1 \block_mem_reg[11][1]  ( .D(n1724), .CLK(clk), .Q(core_block[641])
         );
  DFFPOSX1 \block_mem_reg[11][0]  ( .D(n1723), .CLK(clk), .Q(core_block[640])
         );
  DFFPOSX1 \block_mem_reg[12][31]  ( .D(n1722), .CLK(clk), .Q(core_block[639])
         );
  DFFPOSX1 \block_mem_reg[12][30]  ( .D(n1721), .CLK(clk), .Q(core_block[638])
         );
  DFFPOSX1 \block_mem_reg[12][29]  ( .D(n1720), .CLK(clk), .Q(core_block[637])
         );
  DFFPOSX1 \block_mem_reg[12][28]  ( .D(n1719), .CLK(clk), .Q(core_block[636])
         );
  DFFPOSX1 \block_mem_reg[12][27]  ( .D(n1718), .CLK(clk), .Q(core_block[635])
         );
  DFFPOSX1 \block_mem_reg[12][26]  ( .D(n1717), .CLK(clk), .Q(core_block[634])
         );
  DFFPOSX1 \block_mem_reg[12][25]  ( .D(n1716), .CLK(clk), .Q(core_block[633])
         );
  DFFPOSX1 \block_mem_reg[12][24]  ( .D(n1715), .CLK(clk), .Q(core_block[632])
         );
  DFFPOSX1 \block_mem_reg[12][23]  ( .D(n1714), .CLK(clk), .Q(core_block[631])
         );
  DFFPOSX1 \block_mem_reg[12][22]  ( .D(n1713), .CLK(clk), .Q(core_block[630])
         );
  DFFPOSX1 \block_mem_reg[12][21]  ( .D(n1712), .CLK(clk), .Q(core_block[629])
         );
  DFFPOSX1 \block_mem_reg[12][20]  ( .D(n1711), .CLK(clk), .Q(core_block[628])
         );
  DFFPOSX1 \block_mem_reg[12][19]  ( .D(n1710), .CLK(clk), .Q(core_block[627])
         );
  DFFPOSX1 \block_mem_reg[12][18]  ( .D(n1709), .CLK(clk), .Q(core_block[626])
         );
  DFFPOSX1 \block_mem_reg[12][17]  ( .D(n1708), .CLK(clk), .Q(core_block[625])
         );
  DFFPOSX1 \block_mem_reg[12][16]  ( .D(n1707), .CLK(clk), .Q(core_block[624])
         );
  DFFPOSX1 \block_mem_reg[12][15]  ( .D(n1706), .CLK(clk), .Q(core_block[623])
         );
  DFFPOSX1 \block_mem_reg[12][14]  ( .D(n1705), .CLK(clk), .Q(core_block[622])
         );
  DFFPOSX1 \block_mem_reg[12][13]  ( .D(n1704), .CLK(clk), .Q(core_block[621])
         );
  DFFPOSX1 \block_mem_reg[12][12]  ( .D(n1703), .CLK(clk), .Q(core_block[620])
         );
  DFFPOSX1 \block_mem_reg[12][11]  ( .D(n1702), .CLK(clk), .Q(core_block[619])
         );
  DFFPOSX1 \block_mem_reg[12][10]  ( .D(n1701), .CLK(clk), .Q(core_block[618])
         );
  DFFPOSX1 \block_mem_reg[12][9]  ( .D(n1700), .CLK(clk), .Q(core_block[617])
         );
  DFFPOSX1 \block_mem_reg[12][8]  ( .D(n1699), .CLK(clk), .Q(core_block[616])
         );
  DFFPOSX1 \block_mem_reg[12][7]  ( .D(n1698), .CLK(clk), .Q(core_block[615])
         );
  DFFPOSX1 \block_mem_reg[12][6]  ( .D(n1697), .CLK(clk), .Q(core_block[614])
         );
  DFFPOSX1 \block_mem_reg[12][5]  ( .D(n1696), .CLK(clk), .Q(core_block[613])
         );
  DFFPOSX1 \block_mem_reg[12][4]  ( .D(n1695), .CLK(clk), .Q(core_block[612])
         );
  DFFPOSX1 \block_mem_reg[12][3]  ( .D(n1694), .CLK(clk), .Q(core_block[611])
         );
  DFFPOSX1 \block_mem_reg[12][2]  ( .D(n1693), .CLK(clk), .Q(core_block[610])
         );
  DFFPOSX1 \block_mem_reg[12][1]  ( .D(n1692), .CLK(clk), .Q(core_block[609])
         );
  DFFPOSX1 \block_mem_reg[12][0]  ( .D(n1691), .CLK(clk), .Q(core_block[608])
         );
  DFFPOSX1 \block_mem_reg[13][31]  ( .D(n1690), .CLK(clk), .Q(core_block[607])
         );
  DFFPOSX1 \block_mem_reg[13][30]  ( .D(n1689), .CLK(clk), .Q(core_block[606])
         );
  DFFPOSX1 \block_mem_reg[13][29]  ( .D(n1688), .CLK(clk), .Q(core_block[605])
         );
  DFFPOSX1 \block_mem_reg[13][28]  ( .D(n1687), .CLK(clk), .Q(core_block[604])
         );
  DFFPOSX1 \block_mem_reg[13][27]  ( .D(n1686), .CLK(clk), .Q(core_block[603])
         );
  DFFPOSX1 \block_mem_reg[13][26]  ( .D(n1685), .CLK(clk), .Q(core_block[602])
         );
  DFFPOSX1 \block_mem_reg[13][25]  ( .D(n1684), .CLK(clk), .Q(core_block[601])
         );
  DFFPOSX1 \block_mem_reg[13][24]  ( .D(n1683), .CLK(clk), .Q(core_block[600])
         );
  DFFPOSX1 \block_mem_reg[13][23]  ( .D(n1682), .CLK(clk), .Q(core_block[599])
         );
  DFFPOSX1 \block_mem_reg[13][22]  ( .D(n1681), .CLK(clk), .Q(core_block[598])
         );
  DFFPOSX1 \block_mem_reg[13][21]  ( .D(n1680), .CLK(clk), .Q(core_block[597])
         );
  DFFPOSX1 \block_mem_reg[13][20]  ( .D(n1679), .CLK(clk), .Q(core_block[596])
         );
  DFFPOSX1 \block_mem_reg[13][19]  ( .D(n1678), .CLK(clk), .Q(core_block[595])
         );
  DFFPOSX1 \block_mem_reg[13][18]  ( .D(n1677), .CLK(clk), .Q(core_block[594])
         );
  DFFPOSX1 \block_mem_reg[13][17]  ( .D(n1676), .CLK(clk), .Q(core_block[593])
         );
  DFFPOSX1 \block_mem_reg[13][16]  ( .D(n1675), .CLK(clk), .Q(core_block[592])
         );
  DFFPOSX1 \block_mem_reg[13][15]  ( .D(n1674), .CLK(clk), .Q(core_block[591])
         );
  DFFPOSX1 \block_mem_reg[13][14]  ( .D(n1673), .CLK(clk), .Q(core_block[590])
         );
  DFFPOSX1 \block_mem_reg[13][13]  ( .D(n1672), .CLK(clk), .Q(core_block[589])
         );
  DFFPOSX1 \block_mem_reg[13][12]  ( .D(n1671), .CLK(clk), .Q(core_block[588])
         );
  DFFPOSX1 \block_mem_reg[13][11]  ( .D(n1670), .CLK(clk), .Q(core_block[587])
         );
  DFFPOSX1 \block_mem_reg[13][10]  ( .D(n1669), .CLK(clk), .Q(core_block[586])
         );
  DFFPOSX1 \block_mem_reg[13][9]  ( .D(n1668), .CLK(clk), .Q(core_block[585])
         );
  DFFPOSX1 \block_mem_reg[13][8]  ( .D(n1667), .CLK(clk), .Q(core_block[584])
         );
  DFFPOSX1 \block_mem_reg[13][7]  ( .D(n1666), .CLK(clk), .Q(core_block[583])
         );
  DFFPOSX1 \block_mem_reg[13][6]  ( .D(n1665), .CLK(clk), .Q(core_block[582])
         );
  DFFPOSX1 \block_mem_reg[13][5]  ( .D(n1664), .CLK(clk), .Q(core_block[581])
         );
  DFFPOSX1 \block_mem_reg[13][4]  ( .D(n1663), .CLK(clk), .Q(core_block[580])
         );
  DFFPOSX1 \block_mem_reg[13][3]  ( .D(n1662), .CLK(clk), .Q(core_block[579])
         );
  DFFPOSX1 \block_mem_reg[13][2]  ( .D(n1661), .CLK(clk), .Q(core_block[578])
         );
  DFFPOSX1 \block_mem_reg[13][1]  ( .D(n1660), .CLK(clk), .Q(core_block[577])
         );
  DFFPOSX1 \block_mem_reg[13][0]  ( .D(n1659), .CLK(clk), .Q(core_block[576])
         );
  DFFPOSX1 \block_mem_reg[14][31]  ( .D(n1658), .CLK(clk), .Q(core_block[575])
         );
  DFFPOSX1 \block_mem_reg[14][30]  ( .D(n1657), .CLK(clk), .Q(core_block[574])
         );
  DFFPOSX1 \block_mem_reg[14][29]  ( .D(n1656), .CLK(clk), .Q(core_block[573])
         );
  DFFPOSX1 \block_mem_reg[14][28]  ( .D(n1655), .CLK(clk), .Q(core_block[572])
         );
  DFFPOSX1 \block_mem_reg[14][27]  ( .D(n1654), .CLK(clk), .Q(core_block[571])
         );
  DFFPOSX1 \block_mem_reg[14][26]  ( .D(n1653), .CLK(clk), .Q(core_block[570])
         );
  DFFPOSX1 \block_mem_reg[14][25]  ( .D(n1652), .CLK(clk), .Q(core_block[569])
         );
  DFFPOSX1 \block_mem_reg[14][24]  ( .D(n1651), .CLK(clk), .Q(core_block[568])
         );
  DFFPOSX1 \block_mem_reg[14][23]  ( .D(n1650), .CLK(clk), .Q(core_block[567])
         );
  DFFPOSX1 \block_mem_reg[14][22]  ( .D(n1649), .CLK(clk), .Q(core_block[566])
         );
  DFFPOSX1 \block_mem_reg[14][21]  ( .D(n1648), .CLK(clk), .Q(core_block[565])
         );
  DFFPOSX1 \block_mem_reg[14][20]  ( .D(n1647), .CLK(clk), .Q(core_block[564])
         );
  DFFPOSX1 \block_mem_reg[14][19]  ( .D(n1646), .CLK(clk), .Q(core_block[563])
         );
  DFFPOSX1 \block_mem_reg[14][18]  ( .D(n1645), .CLK(clk), .Q(core_block[562])
         );
  DFFPOSX1 \block_mem_reg[14][17]  ( .D(n1644), .CLK(clk), .Q(core_block[561])
         );
  DFFPOSX1 \block_mem_reg[14][16]  ( .D(n1643), .CLK(clk), .Q(core_block[560])
         );
  DFFPOSX1 \block_mem_reg[14][15]  ( .D(n1642), .CLK(clk), .Q(core_block[559])
         );
  DFFPOSX1 \block_mem_reg[14][14]  ( .D(n1641), .CLK(clk), .Q(core_block[558])
         );
  DFFPOSX1 \block_mem_reg[14][13]  ( .D(n1640), .CLK(clk), .Q(core_block[557])
         );
  DFFPOSX1 \block_mem_reg[14][12]  ( .D(n1639), .CLK(clk), .Q(core_block[556])
         );
  DFFPOSX1 \block_mem_reg[14][11]  ( .D(n1638), .CLK(clk), .Q(core_block[555])
         );
  DFFPOSX1 \block_mem_reg[14][10]  ( .D(n1637), .CLK(clk), .Q(core_block[554])
         );
  DFFPOSX1 \block_mem_reg[14][9]  ( .D(n1636), .CLK(clk), .Q(core_block[553])
         );
  DFFPOSX1 \block_mem_reg[14][8]  ( .D(n1635), .CLK(clk), .Q(core_block[552])
         );
  DFFPOSX1 \block_mem_reg[14][7]  ( .D(n1634), .CLK(clk), .Q(core_block[551])
         );
  DFFPOSX1 \block_mem_reg[14][6]  ( .D(n1633), .CLK(clk), .Q(core_block[550])
         );
  DFFPOSX1 \block_mem_reg[14][5]  ( .D(n1632), .CLK(clk), .Q(core_block[549])
         );
  DFFPOSX1 \block_mem_reg[14][4]  ( .D(n1631), .CLK(clk), .Q(core_block[548])
         );
  DFFPOSX1 \block_mem_reg[14][3]  ( .D(n1630), .CLK(clk), .Q(core_block[547])
         );
  DFFPOSX1 \block_mem_reg[14][2]  ( .D(n1629), .CLK(clk), .Q(core_block[546])
         );
  DFFPOSX1 \block_mem_reg[14][1]  ( .D(n1628), .CLK(clk), .Q(core_block[545])
         );
  DFFPOSX1 \block_mem_reg[14][0]  ( .D(n1627), .CLK(clk), .Q(core_block[544])
         );
  DFFPOSX1 \block_mem_reg[15][31]  ( .D(n1626), .CLK(clk), .Q(core_block[543])
         );
  DFFPOSX1 \block_mem_reg[15][30]  ( .D(n1625), .CLK(clk), .Q(core_block[542])
         );
  DFFPOSX1 \block_mem_reg[15][29]  ( .D(n1624), .CLK(clk), .Q(core_block[541])
         );
  DFFPOSX1 \block_mem_reg[15][28]  ( .D(n1623), .CLK(clk), .Q(core_block[540])
         );
  DFFPOSX1 \block_mem_reg[15][27]  ( .D(n1622), .CLK(clk), .Q(core_block[539])
         );
  DFFPOSX1 \block_mem_reg[15][26]  ( .D(n1621), .CLK(clk), .Q(core_block[538])
         );
  DFFPOSX1 \block_mem_reg[15][25]  ( .D(n1620), .CLK(clk), .Q(core_block[537])
         );
  DFFPOSX1 \block_mem_reg[15][24]  ( .D(n1619), .CLK(clk), .Q(core_block[536])
         );
  DFFPOSX1 \block_mem_reg[15][23]  ( .D(n1618), .CLK(clk), .Q(core_block[535])
         );
  DFFPOSX1 \block_mem_reg[15][22]  ( .D(n1617), .CLK(clk), .Q(core_block[534])
         );
  DFFPOSX1 \block_mem_reg[15][21]  ( .D(n1616), .CLK(clk), .Q(core_block[533])
         );
  DFFPOSX1 \block_mem_reg[15][20]  ( .D(n1615), .CLK(clk), .Q(core_block[532])
         );
  DFFPOSX1 \block_mem_reg[15][19]  ( .D(n1614), .CLK(clk), .Q(core_block[531])
         );
  DFFPOSX1 \block_mem_reg[15][18]  ( .D(n1613), .CLK(clk), .Q(core_block[530])
         );
  DFFPOSX1 \block_mem_reg[15][17]  ( .D(n1612), .CLK(clk), .Q(core_block[529])
         );
  DFFPOSX1 \block_mem_reg[15][16]  ( .D(n1611), .CLK(clk), .Q(core_block[528])
         );
  DFFPOSX1 \block_mem_reg[15][15]  ( .D(n1610), .CLK(clk), .Q(core_block[527])
         );
  DFFPOSX1 \block_mem_reg[15][14]  ( .D(n1609), .CLK(clk), .Q(core_block[526])
         );
  DFFPOSX1 \block_mem_reg[15][13]  ( .D(n1608), .CLK(clk), .Q(core_block[525])
         );
  DFFPOSX1 \block_mem_reg[15][12]  ( .D(n1607), .CLK(clk), .Q(core_block[524])
         );
  DFFPOSX1 \block_mem_reg[15][11]  ( .D(n1606), .CLK(clk), .Q(core_block[523])
         );
  DFFPOSX1 \block_mem_reg[15][10]  ( .D(n1605), .CLK(clk), .Q(core_block[522])
         );
  DFFPOSX1 \block_mem_reg[15][9]  ( .D(n1604), .CLK(clk), .Q(core_block[521])
         );
  DFFPOSX1 \block_mem_reg[15][8]  ( .D(n1603), .CLK(clk), .Q(core_block[520])
         );
  DFFPOSX1 \block_mem_reg[15][7]  ( .D(n1602), .CLK(clk), .Q(core_block[519])
         );
  DFFPOSX1 \block_mem_reg[15][6]  ( .D(n1601), .CLK(clk), .Q(core_block[518])
         );
  DFFPOSX1 \block_mem_reg[15][5]  ( .D(n1600), .CLK(clk), .Q(core_block[517])
         );
  DFFPOSX1 \block_mem_reg[15][4]  ( .D(n1599), .CLK(clk), .Q(core_block[516])
         );
  DFFPOSX1 \block_mem_reg[15][3]  ( .D(n1598), .CLK(clk), .Q(core_block[515])
         );
  DFFPOSX1 \block_mem_reg[15][2]  ( .D(n1597), .CLK(clk), .Q(core_block[514])
         );
  DFFPOSX1 \block_mem_reg[15][1]  ( .D(n1596), .CLK(clk), .Q(core_block[513])
         );
  DFFPOSX1 \block_mem_reg[15][0]  ( .D(n1595), .CLK(clk), .Q(core_block[512])
         );
  DFFPOSX1 \block_mem_reg[16][31]  ( .D(n1594), .CLK(clk), .Q(core_block[511])
         );
  DFFPOSX1 \block_mem_reg[16][30]  ( .D(n1593), .CLK(clk), .Q(core_block[510])
         );
  DFFPOSX1 \block_mem_reg[16][29]  ( .D(n1592), .CLK(clk), .Q(core_block[509])
         );
  DFFPOSX1 \block_mem_reg[16][28]  ( .D(n1591), .CLK(clk), .Q(core_block[508])
         );
  DFFPOSX1 \block_mem_reg[16][27]  ( .D(n1590), .CLK(clk), .Q(core_block[507])
         );
  DFFPOSX1 \block_mem_reg[16][26]  ( .D(n1589), .CLK(clk), .Q(core_block[506])
         );
  DFFPOSX1 \block_mem_reg[16][25]  ( .D(n1588), .CLK(clk), .Q(core_block[505])
         );
  DFFPOSX1 \block_mem_reg[16][24]  ( .D(n1587), .CLK(clk), .Q(core_block[504])
         );
  DFFPOSX1 \block_mem_reg[16][23]  ( .D(n1586), .CLK(clk), .Q(core_block[503])
         );
  DFFPOSX1 \block_mem_reg[16][22]  ( .D(n1585), .CLK(clk), .Q(core_block[502])
         );
  DFFPOSX1 \block_mem_reg[16][21]  ( .D(n1584), .CLK(clk), .Q(core_block[501])
         );
  DFFPOSX1 \block_mem_reg[16][20]  ( .D(n1583), .CLK(clk), .Q(core_block[500])
         );
  DFFPOSX1 \block_mem_reg[16][19]  ( .D(n1582), .CLK(clk), .Q(core_block[499])
         );
  DFFPOSX1 \block_mem_reg[16][18]  ( .D(n1581), .CLK(clk), .Q(core_block[498])
         );
  DFFPOSX1 \block_mem_reg[16][17]  ( .D(n1580), .CLK(clk), .Q(core_block[497])
         );
  DFFPOSX1 \block_mem_reg[16][16]  ( .D(n1579), .CLK(clk), .Q(core_block[496])
         );
  DFFPOSX1 \block_mem_reg[16][15]  ( .D(n1578), .CLK(clk), .Q(core_block[495])
         );
  DFFPOSX1 \block_mem_reg[16][14]  ( .D(n1577), .CLK(clk), .Q(core_block[494])
         );
  DFFPOSX1 \block_mem_reg[16][13]  ( .D(n1576), .CLK(clk), .Q(core_block[493])
         );
  DFFPOSX1 \block_mem_reg[16][12]  ( .D(n1575), .CLK(clk), .Q(core_block[492])
         );
  DFFPOSX1 \block_mem_reg[16][11]  ( .D(n1574), .CLK(clk), .Q(core_block[491])
         );
  DFFPOSX1 \block_mem_reg[16][10]  ( .D(n1573), .CLK(clk), .Q(core_block[490])
         );
  DFFPOSX1 \block_mem_reg[16][9]  ( .D(n1572), .CLK(clk), .Q(core_block[489])
         );
  DFFPOSX1 \block_mem_reg[16][8]  ( .D(n1571), .CLK(clk), .Q(core_block[488])
         );
  DFFPOSX1 \block_mem_reg[16][7]  ( .D(n1570), .CLK(clk), .Q(core_block[487])
         );
  DFFPOSX1 \block_mem_reg[16][6]  ( .D(n1569), .CLK(clk), .Q(core_block[486])
         );
  DFFPOSX1 \block_mem_reg[16][5]  ( .D(n1568), .CLK(clk), .Q(core_block[485])
         );
  DFFPOSX1 \block_mem_reg[16][4]  ( .D(n1567), .CLK(clk), .Q(core_block[484])
         );
  DFFPOSX1 \block_mem_reg[16][3]  ( .D(n1566), .CLK(clk), .Q(core_block[483])
         );
  DFFPOSX1 \block_mem_reg[16][2]  ( .D(n1565), .CLK(clk), .Q(core_block[482])
         );
  DFFPOSX1 \block_mem_reg[16][1]  ( .D(n1564), .CLK(clk), .Q(core_block[481])
         );
  DFFPOSX1 \block_mem_reg[16][0]  ( .D(n1563), .CLK(clk), .Q(core_block[480])
         );
  DFFPOSX1 \block_mem_reg[17][31]  ( .D(n1562), .CLK(clk), .Q(core_block[479])
         );
  DFFPOSX1 \block_mem_reg[17][30]  ( .D(n1561), .CLK(clk), .Q(core_block[478])
         );
  DFFPOSX1 \block_mem_reg[17][29]  ( .D(n1560), .CLK(clk), .Q(core_block[477])
         );
  DFFPOSX1 \block_mem_reg[17][28]  ( .D(n1559), .CLK(clk), .Q(core_block[476])
         );
  DFFPOSX1 \block_mem_reg[17][27]  ( .D(n1558), .CLK(clk), .Q(core_block[475])
         );
  DFFPOSX1 \block_mem_reg[17][26]  ( .D(n1557), .CLK(clk), .Q(core_block[474])
         );
  DFFPOSX1 \block_mem_reg[17][25]  ( .D(n1556), .CLK(clk), .Q(core_block[473])
         );
  DFFPOSX1 \block_mem_reg[17][24]  ( .D(n1555), .CLK(clk), .Q(core_block[472])
         );
  DFFPOSX1 \block_mem_reg[17][23]  ( .D(n1554), .CLK(clk), .Q(core_block[471])
         );
  DFFPOSX1 \block_mem_reg[17][22]  ( .D(n1553), .CLK(clk), .Q(core_block[470])
         );
  DFFPOSX1 \block_mem_reg[17][21]  ( .D(n1552), .CLK(clk), .Q(core_block[469])
         );
  DFFPOSX1 \block_mem_reg[17][20]  ( .D(n1551), .CLK(clk), .Q(core_block[468])
         );
  DFFPOSX1 \block_mem_reg[17][19]  ( .D(n1550), .CLK(clk), .Q(core_block[467])
         );
  DFFPOSX1 \block_mem_reg[17][18]  ( .D(n1549), .CLK(clk), .Q(core_block[466])
         );
  DFFPOSX1 \block_mem_reg[17][17]  ( .D(n1548), .CLK(clk), .Q(core_block[465])
         );
  DFFPOSX1 \block_mem_reg[17][16]  ( .D(n1547), .CLK(clk), .Q(core_block[464])
         );
  DFFPOSX1 \block_mem_reg[17][15]  ( .D(n1546), .CLK(clk), .Q(core_block[463])
         );
  DFFPOSX1 \block_mem_reg[17][14]  ( .D(n1545), .CLK(clk), .Q(core_block[462])
         );
  DFFPOSX1 \block_mem_reg[17][13]  ( .D(n1544), .CLK(clk), .Q(core_block[461])
         );
  DFFPOSX1 \block_mem_reg[17][12]  ( .D(n1543), .CLK(clk), .Q(core_block[460])
         );
  DFFPOSX1 \block_mem_reg[17][11]  ( .D(n1542), .CLK(clk), .Q(core_block[459])
         );
  DFFPOSX1 \block_mem_reg[17][10]  ( .D(n1541), .CLK(clk), .Q(core_block[458])
         );
  DFFPOSX1 \block_mem_reg[17][9]  ( .D(n1540), .CLK(clk), .Q(core_block[457])
         );
  DFFPOSX1 \block_mem_reg[17][8]  ( .D(n1539), .CLK(clk), .Q(core_block[456])
         );
  DFFPOSX1 \block_mem_reg[17][7]  ( .D(n1538), .CLK(clk), .Q(core_block[455])
         );
  DFFPOSX1 \block_mem_reg[17][6]  ( .D(n1537), .CLK(clk), .Q(core_block[454])
         );
  DFFPOSX1 \block_mem_reg[17][5]  ( .D(n1536), .CLK(clk), .Q(core_block[453])
         );
  DFFPOSX1 \block_mem_reg[17][4]  ( .D(n1535), .CLK(clk), .Q(core_block[452])
         );
  DFFPOSX1 \block_mem_reg[17][3]  ( .D(n1534), .CLK(clk), .Q(core_block[451])
         );
  DFFPOSX1 \block_mem_reg[17][2]  ( .D(n1533), .CLK(clk), .Q(core_block[450])
         );
  DFFPOSX1 \block_mem_reg[17][1]  ( .D(n1532), .CLK(clk), .Q(core_block[449])
         );
  DFFPOSX1 \block_mem_reg[17][0]  ( .D(n1531), .CLK(clk), .Q(core_block[448])
         );
  DFFPOSX1 \block_mem_reg[18][31]  ( .D(n1530), .CLK(clk), .Q(core_block[447])
         );
  DFFPOSX1 \block_mem_reg[18][30]  ( .D(n1529), .CLK(clk), .Q(core_block[446])
         );
  DFFPOSX1 \block_mem_reg[18][29]  ( .D(n1528), .CLK(clk), .Q(core_block[445])
         );
  DFFPOSX1 \block_mem_reg[18][28]  ( .D(n1527), .CLK(clk), .Q(core_block[444])
         );
  DFFPOSX1 \block_mem_reg[18][27]  ( .D(n1526), .CLK(clk), .Q(core_block[443])
         );
  DFFPOSX1 \block_mem_reg[18][26]  ( .D(n1525), .CLK(clk), .Q(core_block[442])
         );
  DFFPOSX1 \block_mem_reg[18][25]  ( .D(n1524), .CLK(clk), .Q(core_block[441])
         );
  DFFPOSX1 \block_mem_reg[18][24]  ( .D(n1523), .CLK(clk), .Q(core_block[440])
         );
  DFFPOSX1 \block_mem_reg[18][23]  ( .D(n1522), .CLK(clk), .Q(core_block[439])
         );
  DFFPOSX1 \block_mem_reg[18][22]  ( .D(n1521), .CLK(clk), .Q(core_block[438])
         );
  DFFPOSX1 \block_mem_reg[18][21]  ( .D(n1520), .CLK(clk), .Q(core_block[437])
         );
  DFFPOSX1 \block_mem_reg[18][20]  ( .D(n1519), .CLK(clk), .Q(core_block[436])
         );
  DFFPOSX1 \block_mem_reg[18][19]  ( .D(n1518), .CLK(clk), .Q(core_block[435])
         );
  DFFPOSX1 \block_mem_reg[18][18]  ( .D(n1517), .CLK(clk), .Q(core_block[434])
         );
  DFFPOSX1 \block_mem_reg[18][17]  ( .D(n1516), .CLK(clk), .Q(core_block[433])
         );
  DFFPOSX1 \block_mem_reg[18][16]  ( .D(n1515), .CLK(clk), .Q(core_block[432])
         );
  DFFPOSX1 \block_mem_reg[18][15]  ( .D(n1514), .CLK(clk), .Q(core_block[431])
         );
  DFFPOSX1 \block_mem_reg[18][14]  ( .D(n1513), .CLK(clk), .Q(core_block[430])
         );
  DFFPOSX1 \block_mem_reg[18][13]  ( .D(n1512), .CLK(clk), .Q(core_block[429])
         );
  DFFPOSX1 \block_mem_reg[18][12]  ( .D(n1511), .CLK(clk), .Q(core_block[428])
         );
  DFFPOSX1 \block_mem_reg[18][11]  ( .D(n1510), .CLK(clk), .Q(core_block[427])
         );
  DFFPOSX1 \block_mem_reg[18][10]  ( .D(n1509), .CLK(clk), .Q(core_block[426])
         );
  DFFPOSX1 \block_mem_reg[18][9]  ( .D(n1508), .CLK(clk), .Q(core_block[425])
         );
  DFFPOSX1 \block_mem_reg[18][8]  ( .D(n1507), .CLK(clk), .Q(core_block[424])
         );
  DFFPOSX1 \block_mem_reg[18][7]  ( .D(n1506), .CLK(clk), .Q(core_block[423])
         );
  DFFPOSX1 \block_mem_reg[18][6]  ( .D(n1505), .CLK(clk), .Q(core_block[422])
         );
  DFFPOSX1 \block_mem_reg[18][5]  ( .D(n1504), .CLK(clk), .Q(core_block[421])
         );
  DFFPOSX1 \block_mem_reg[18][4]  ( .D(n1503), .CLK(clk), .Q(core_block[420])
         );
  DFFPOSX1 \block_mem_reg[18][3]  ( .D(n1502), .CLK(clk), .Q(core_block[419])
         );
  DFFPOSX1 \block_mem_reg[18][2]  ( .D(n1501), .CLK(clk), .Q(core_block[418])
         );
  DFFPOSX1 \block_mem_reg[18][1]  ( .D(n1500), .CLK(clk), .Q(core_block[417])
         );
  DFFPOSX1 \block_mem_reg[18][0]  ( .D(n1499), .CLK(clk), .Q(core_block[416])
         );
  DFFPOSX1 \block_mem_reg[19][31]  ( .D(n1498), .CLK(clk), .Q(core_block[415])
         );
  DFFPOSX1 \block_mem_reg[19][30]  ( .D(n1497), .CLK(clk), .Q(core_block[414])
         );
  DFFPOSX1 \block_mem_reg[19][29]  ( .D(n1496), .CLK(clk), .Q(core_block[413])
         );
  DFFPOSX1 \block_mem_reg[19][28]  ( .D(n1495), .CLK(clk), .Q(core_block[412])
         );
  DFFPOSX1 \block_mem_reg[19][27]  ( .D(n1494), .CLK(clk), .Q(core_block[411])
         );
  DFFPOSX1 \block_mem_reg[19][26]  ( .D(n1493), .CLK(clk), .Q(core_block[410])
         );
  DFFPOSX1 \block_mem_reg[19][25]  ( .D(n1492), .CLK(clk), .Q(core_block[409])
         );
  DFFPOSX1 \block_mem_reg[19][24]  ( .D(n1491), .CLK(clk), .Q(core_block[408])
         );
  DFFPOSX1 \block_mem_reg[19][23]  ( .D(n1490), .CLK(clk), .Q(core_block[407])
         );
  DFFPOSX1 \block_mem_reg[19][22]  ( .D(n1489), .CLK(clk), .Q(core_block[406])
         );
  DFFPOSX1 \block_mem_reg[19][21]  ( .D(n1488), .CLK(clk), .Q(core_block[405])
         );
  DFFPOSX1 \block_mem_reg[19][20]  ( .D(n1487), .CLK(clk), .Q(core_block[404])
         );
  DFFPOSX1 \block_mem_reg[19][19]  ( .D(n1486), .CLK(clk), .Q(core_block[403])
         );
  DFFPOSX1 \block_mem_reg[19][18]  ( .D(n1485), .CLK(clk), .Q(core_block[402])
         );
  DFFPOSX1 \block_mem_reg[19][17]  ( .D(n1484), .CLK(clk), .Q(core_block[401])
         );
  DFFPOSX1 \block_mem_reg[19][16]  ( .D(n1483), .CLK(clk), .Q(core_block[400])
         );
  DFFPOSX1 \block_mem_reg[19][15]  ( .D(n1482), .CLK(clk), .Q(core_block[399])
         );
  DFFPOSX1 \block_mem_reg[19][14]  ( .D(n1481), .CLK(clk), .Q(core_block[398])
         );
  DFFPOSX1 \block_mem_reg[19][13]  ( .D(n1480), .CLK(clk), .Q(core_block[397])
         );
  DFFPOSX1 \block_mem_reg[19][12]  ( .D(n1479), .CLK(clk), .Q(core_block[396])
         );
  DFFPOSX1 \block_mem_reg[19][11]  ( .D(n1478), .CLK(clk), .Q(core_block[395])
         );
  DFFPOSX1 \block_mem_reg[19][10]  ( .D(n1477), .CLK(clk), .Q(core_block[394])
         );
  DFFPOSX1 \block_mem_reg[19][9]  ( .D(n1476), .CLK(clk), .Q(core_block[393])
         );
  DFFPOSX1 \block_mem_reg[19][8]  ( .D(n1475), .CLK(clk), .Q(core_block[392])
         );
  DFFPOSX1 \block_mem_reg[19][7]  ( .D(n1474), .CLK(clk), .Q(core_block[391])
         );
  DFFPOSX1 \block_mem_reg[19][6]  ( .D(n1473), .CLK(clk), .Q(core_block[390])
         );
  DFFPOSX1 \block_mem_reg[19][5]  ( .D(n1472), .CLK(clk), .Q(core_block[389])
         );
  DFFPOSX1 \block_mem_reg[19][4]  ( .D(n1471), .CLK(clk), .Q(core_block[388])
         );
  DFFPOSX1 \block_mem_reg[19][3]  ( .D(n1470), .CLK(clk), .Q(core_block[387])
         );
  DFFPOSX1 \block_mem_reg[19][2]  ( .D(n1469), .CLK(clk), .Q(core_block[386])
         );
  DFFPOSX1 \block_mem_reg[19][1]  ( .D(n1468), .CLK(clk), .Q(core_block[385])
         );
  DFFPOSX1 \block_mem_reg[19][0]  ( .D(n1467), .CLK(clk), .Q(core_block[384])
         );
  DFFPOSX1 \block_mem_reg[20][31]  ( .D(n1466), .CLK(clk), .Q(core_block[383])
         );
  DFFPOSX1 \block_mem_reg[20][30]  ( .D(n1465), .CLK(clk), .Q(core_block[382])
         );
  DFFPOSX1 \block_mem_reg[20][29]  ( .D(n1464), .CLK(clk), .Q(core_block[381])
         );
  DFFPOSX1 \block_mem_reg[20][28]  ( .D(n1463), .CLK(clk), .Q(core_block[380])
         );
  DFFPOSX1 \block_mem_reg[20][27]  ( .D(n1462), .CLK(clk), .Q(core_block[379])
         );
  DFFPOSX1 \block_mem_reg[20][26]  ( .D(n1461), .CLK(clk), .Q(core_block[378])
         );
  DFFPOSX1 \block_mem_reg[20][25]  ( .D(n1460), .CLK(clk), .Q(core_block[377])
         );
  DFFPOSX1 \block_mem_reg[20][24]  ( .D(n1459), .CLK(clk), .Q(core_block[376])
         );
  DFFPOSX1 \block_mem_reg[20][23]  ( .D(n1458), .CLK(clk), .Q(core_block[375])
         );
  DFFPOSX1 \block_mem_reg[20][22]  ( .D(n1457), .CLK(clk), .Q(core_block[374])
         );
  DFFPOSX1 \block_mem_reg[20][21]  ( .D(n1456), .CLK(clk), .Q(core_block[373])
         );
  DFFPOSX1 \block_mem_reg[20][20]  ( .D(n1455), .CLK(clk), .Q(core_block[372])
         );
  DFFPOSX1 \block_mem_reg[20][19]  ( .D(n1454), .CLK(clk), .Q(core_block[371])
         );
  DFFPOSX1 \block_mem_reg[20][18]  ( .D(n1453), .CLK(clk), .Q(core_block[370])
         );
  DFFPOSX1 \block_mem_reg[20][17]  ( .D(n1452), .CLK(clk), .Q(core_block[369])
         );
  DFFPOSX1 \block_mem_reg[20][16]  ( .D(n1451), .CLK(clk), .Q(core_block[368])
         );
  DFFPOSX1 \block_mem_reg[20][15]  ( .D(n1450), .CLK(clk), .Q(core_block[367])
         );
  DFFPOSX1 \block_mem_reg[20][14]  ( .D(n1449), .CLK(clk), .Q(core_block[366])
         );
  DFFPOSX1 \block_mem_reg[20][13]  ( .D(n1448), .CLK(clk), .Q(core_block[365])
         );
  DFFPOSX1 \block_mem_reg[20][12]  ( .D(n1447), .CLK(clk), .Q(core_block[364])
         );
  DFFPOSX1 \block_mem_reg[20][11]  ( .D(n1446), .CLK(clk), .Q(core_block[363])
         );
  DFFPOSX1 \block_mem_reg[20][10]  ( .D(n1445), .CLK(clk), .Q(core_block[362])
         );
  DFFPOSX1 \block_mem_reg[20][9]  ( .D(n1444), .CLK(clk), .Q(core_block[361])
         );
  DFFPOSX1 \block_mem_reg[20][8]  ( .D(n1443), .CLK(clk), .Q(core_block[360])
         );
  DFFPOSX1 \block_mem_reg[20][7]  ( .D(n1442), .CLK(clk), .Q(core_block[359])
         );
  DFFPOSX1 \block_mem_reg[20][6]  ( .D(n1441), .CLK(clk), .Q(core_block[358])
         );
  DFFPOSX1 \block_mem_reg[20][5]  ( .D(n1440), .CLK(clk), .Q(core_block[357])
         );
  DFFPOSX1 \block_mem_reg[20][4]  ( .D(n1439), .CLK(clk), .Q(core_block[356])
         );
  DFFPOSX1 \block_mem_reg[20][3]  ( .D(n1438), .CLK(clk), .Q(core_block[355])
         );
  DFFPOSX1 \block_mem_reg[20][2]  ( .D(n1437), .CLK(clk), .Q(core_block[354])
         );
  DFFPOSX1 \block_mem_reg[20][1]  ( .D(n1436), .CLK(clk), .Q(core_block[353])
         );
  DFFPOSX1 \block_mem_reg[20][0]  ( .D(n1435), .CLK(clk), .Q(core_block[352])
         );
  DFFPOSX1 \block_mem_reg[21][31]  ( .D(n1434), .CLK(clk), .Q(core_block[351])
         );
  DFFPOSX1 \block_mem_reg[21][30]  ( .D(n1433), .CLK(clk), .Q(core_block[350])
         );
  DFFPOSX1 \block_mem_reg[21][29]  ( .D(n1432), .CLK(clk), .Q(core_block[349])
         );
  DFFPOSX1 \block_mem_reg[21][28]  ( .D(n1431), .CLK(clk), .Q(core_block[348])
         );
  DFFPOSX1 \block_mem_reg[21][27]  ( .D(n1430), .CLK(clk), .Q(core_block[347])
         );
  DFFPOSX1 \block_mem_reg[21][26]  ( .D(n1429), .CLK(clk), .Q(core_block[346])
         );
  DFFPOSX1 \block_mem_reg[21][25]  ( .D(n1428), .CLK(clk), .Q(core_block[345])
         );
  DFFPOSX1 \block_mem_reg[21][24]  ( .D(n1427), .CLK(clk), .Q(core_block[344])
         );
  DFFPOSX1 \block_mem_reg[21][23]  ( .D(n1426), .CLK(clk), .Q(core_block[343])
         );
  DFFPOSX1 \block_mem_reg[21][22]  ( .D(n1425), .CLK(clk), .Q(core_block[342])
         );
  DFFPOSX1 \block_mem_reg[21][21]  ( .D(n1424), .CLK(clk), .Q(core_block[341])
         );
  DFFPOSX1 \block_mem_reg[21][20]  ( .D(n1423), .CLK(clk), .Q(core_block[340])
         );
  DFFPOSX1 \block_mem_reg[21][19]  ( .D(n1422), .CLK(clk), .Q(core_block[339])
         );
  DFFPOSX1 \block_mem_reg[21][18]  ( .D(n1421), .CLK(clk), .Q(core_block[338])
         );
  DFFPOSX1 \block_mem_reg[21][17]  ( .D(n1420), .CLK(clk), .Q(core_block[337])
         );
  DFFPOSX1 \block_mem_reg[21][16]  ( .D(n1419), .CLK(clk), .Q(core_block[336])
         );
  DFFPOSX1 \block_mem_reg[21][15]  ( .D(n1418), .CLK(clk), .Q(core_block[335])
         );
  DFFPOSX1 \block_mem_reg[21][14]  ( .D(n1417), .CLK(clk), .Q(core_block[334])
         );
  DFFPOSX1 \block_mem_reg[21][13]  ( .D(n1416), .CLK(clk), .Q(core_block[333])
         );
  DFFPOSX1 \block_mem_reg[21][12]  ( .D(n1415), .CLK(clk), .Q(core_block[332])
         );
  DFFPOSX1 \block_mem_reg[21][11]  ( .D(n1414), .CLK(clk), .Q(core_block[331])
         );
  DFFPOSX1 \block_mem_reg[21][10]  ( .D(n1413), .CLK(clk), .Q(core_block[330])
         );
  DFFPOSX1 \block_mem_reg[21][9]  ( .D(n1412), .CLK(clk), .Q(core_block[329])
         );
  DFFPOSX1 \block_mem_reg[21][8]  ( .D(n1411), .CLK(clk), .Q(core_block[328])
         );
  DFFPOSX1 \block_mem_reg[21][7]  ( .D(n1410), .CLK(clk), .Q(core_block[327])
         );
  DFFPOSX1 \block_mem_reg[21][6]  ( .D(n1409), .CLK(clk), .Q(core_block[326])
         );
  DFFPOSX1 \block_mem_reg[21][5]  ( .D(n1408), .CLK(clk), .Q(core_block[325])
         );
  DFFPOSX1 \block_mem_reg[21][4]  ( .D(n1407), .CLK(clk), .Q(core_block[324])
         );
  DFFPOSX1 \block_mem_reg[21][3]  ( .D(n1406), .CLK(clk), .Q(core_block[323])
         );
  DFFPOSX1 \block_mem_reg[21][2]  ( .D(n1405), .CLK(clk), .Q(core_block[322])
         );
  DFFPOSX1 \block_mem_reg[21][1]  ( .D(n1404), .CLK(clk), .Q(core_block[321])
         );
  DFFPOSX1 \block_mem_reg[21][0]  ( .D(n1403), .CLK(clk), .Q(core_block[320])
         );
  DFFPOSX1 \block_mem_reg[22][31]  ( .D(n1402), .CLK(clk), .Q(core_block[319])
         );
  DFFPOSX1 \block_mem_reg[22][30]  ( .D(n1401), .CLK(clk), .Q(core_block[318])
         );
  DFFPOSX1 \block_mem_reg[22][29]  ( .D(n1400), .CLK(clk), .Q(core_block[317])
         );
  DFFPOSX1 \block_mem_reg[22][28]  ( .D(n1399), .CLK(clk), .Q(core_block[316])
         );
  DFFPOSX1 \block_mem_reg[22][27]  ( .D(n1398), .CLK(clk), .Q(core_block[315])
         );
  DFFPOSX1 \block_mem_reg[22][26]  ( .D(n1397), .CLK(clk), .Q(core_block[314])
         );
  DFFPOSX1 \block_mem_reg[22][25]  ( .D(n1396), .CLK(clk), .Q(core_block[313])
         );
  DFFPOSX1 \block_mem_reg[22][24]  ( .D(n1395), .CLK(clk), .Q(core_block[312])
         );
  DFFPOSX1 \block_mem_reg[22][23]  ( .D(n1394), .CLK(clk), .Q(core_block[311])
         );
  DFFPOSX1 \block_mem_reg[22][22]  ( .D(n1393), .CLK(clk), .Q(core_block[310])
         );
  DFFPOSX1 \block_mem_reg[22][21]  ( .D(n1392), .CLK(clk), .Q(core_block[309])
         );
  DFFPOSX1 \block_mem_reg[22][20]  ( .D(n1391), .CLK(clk), .Q(core_block[308])
         );
  DFFPOSX1 \block_mem_reg[22][19]  ( .D(n1390), .CLK(clk), .Q(core_block[307])
         );
  DFFPOSX1 \block_mem_reg[22][18]  ( .D(n1389), .CLK(clk), .Q(core_block[306])
         );
  DFFPOSX1 \block_mem_reg[22][17]  ( .D(n1388), .CLK(clk), .Q(core_block[305])
         );
  DFFPOSX1 \block_mem_reg[22][16]  ( .D(n1387), .CLK(clk), .Q(core_block[304])
         );
  DFFPOSX1 \block_mem_reg[22][15]  ( .D(n1386), .CLK(clk), .Q(core_block[303])
         );
  DFFPOSX1 \block_mem_reg[22][14]  ( .D(n1385), .CLK(clk), .Q(core_block[302])
         );
  DFFPOSX1 \block_mem_reg[22][13]  ( .D(n1384), .CLK(clk), .Q(core_block[301])
         );
  DFFPOSX1 \block_mem_reg[22][12]  ( .D(n1383), .CLK(clk), .Q(core_block[300])
         );
  DFFPOSX1 \block_mem_reg[22][11]  ( .D(n1382), .CLK(clk), .Q(core_block[299])
         );
  DFFPOSX1 \block_mem_reg[22][10]  ( .D(n1381), .CLK(clk), .Q(core_block[298])
         );
  DFFPOSX1 \block_mem_reg[22][9]  ( .D(n1380), .CLK(clk), .Q(core_block[297])
         );
  DFFPOSX1 \block_mem_reg[22][8]  ( .D(n1379), .CLK(clk), .Q(core_block[296])
         );
  DFFPOSX1 \block_mem_reg[22][7]  ( .D(n1378), .CLK(clk), .Q(core_block[295])
         );
  DFFPOSX1 \block_mem_reg[22][6]  ( .D(n1377), .CLK(clk), .Q(core_block[294])
         );
  DFFPOSX1 \block_mem_reg[22][5]  ( .D(n1376), .CLK(clk), .Q(core_block[293])
         );
  DFFPOSX1 \block_mem_reg[22][4]  ( .D(n1375), .CLK(clk), .Q(core_block[292])
         );
  DFFPOSX1 \block_mem_reg[22][3]  ( .D(n1374), .CLK(clk), .Q(core_block[291])
         );
  DFFPOSX1 \block_mem_reg[22][2]  ( .D(n1373), .CLK(clk), .Q(core_block[290])
         );
  DFFPOSX1 \block_mem_reg[22][1]  ( .D(n1372), .CLK(clk), .Q(core_block[289])
         );
  DFFPOSX1 \block_mem_reg[22][0]  ( .D(n1371), .CLK(clk), .Q(core_block[288])
         );
  DFFPOSX1 \block_mem_reg[23][31]  ( .D(n1370), .CLK(clk), .Q(core_block[287])
         );
  DFFPOSX1 \block_mem_reg[23][30]  ( .D(n1369), .CLK(clk), .Q(core_block[286])
         );
  DFFPOSX1 \block_mem_reg[23][29]  ( .D(n1368), .CLK(clk), .Q(core_block[285])
         );
  DFFPOSX1 \block_mem_reg[23][28]  ( .D(n1367), .CLK(clk), .Q(core_block[284])
         );
  DFFPOSX1 \block_mem_reg[23][27]  ( .D(n1366), .CLK(clk), .Q(core_block[283])
         );
  DFFPOSX1 \block_mem_reg[23][26]  ( .D(n1365), .CLK(clk), .Q(core_block[282])
         );
  DFFPOSX1 \block_mem_reg[23][25]  ( .D(n1364), .CLK(clk), .Q(core_block[281])
         );
  DFFPOSX1 \block_mem_reg[23][24]  ( .D(n1363), .CLK(clk), .Q(core_block[280])
         );
  DFFPOSX1 \block_mem_reg[23][23]  ( .D(n1362), .CLK(clk), .Q(core_block[279])
         );
  DFFPOSX1 \block_mem_reg[23][22]  ( .D(n1361), .CLK(clk), .Q(core_block[278])
         );
  DFFPOSX1 \block_mem_reg[23][21]  ( .D(n1360), .CLK(clk), .Q(core_block[277])
         );
  DFFPOSX1 \block_mem_reg[23][20]  ( .D(n1359), .CLK(clk), .Q(core_block[276])
         );
  DFFPOSX1 \block_mem_reg[23][19]  ( .D(n1358), .CLK(clk), .Q(core_block[275])
         );
  DFFPOSX1 \block_mem_reg[23][18]  ( .D(n1357), .CLK(clk), .Q(core_block[274])
         );
  DFFPOSX1 \block_mem_reg[23][17]  ( .D(n1356), .CLK(clk), .Q(core_block[273])
         );
  DFFPOSX1 \block_mem_reg[23][16]  ( .D(n1355), .CLK(clk), .Q(core_block[272])
         );
  DFFPOSX1 \block_mem_reg[23][15]  ( .D(n1354), .CLK(clk), .Q(core_block[271])
         );
  DFFPOSX1 \block_mem_reg[23][14]  ( .D(n1353), .CLK(clk), .Q(core_block[270])
         );
  DFFPOSX1 \block_mem_reg[23][13]  ( .D(n1352), .CLK(clk), .Q(core_block[269])
         );
  DFFPOSX1 \block_mem_reg[23][12]  ( .D(n1351), .CLK(clk), .Q(core_block[268])
         );
  DFFPOSX1 \block_mem_reg[23][11]  ( .D(n1350), .CLK(clk), .Q(core_block[267])
         );
  DFFPOSX1 \block_mem_reg[23][10]  ( .D(n1349), .CLK(clk), .Q(core_block[266])
         );
  DFFPOSX1 \block_mem_reg[23][9]  ( .D(n1348), .CLK(clk), .Q(core_block[265])
         );
  DFFPOSX1 \block_mem_reg[23][8]  ( .D(n1347), .CLK(clk), .Q(core_block[264])
         );
  DFFPOSX1 \block_mem_reg[23][7]  ( .D(n1346), .CLK(clk), .Q(core_block[263])
         );
  DFFPOSX1 \block_mem_reg[23][6]  ( .D(n1345), .CLK(clk), .Q(core_block[262])
         );
  DFFPOSX1 \block_mem_reg[23][5]  ( .D(n1344), .CLK(clk), .Q(core_block[261])
         );
  DFFPOSX1 \block_mem_reg[23][4]  ( .D(n1343), .CLK(clk), .Q(core_block[260])
         );
  DFFPOSX1 \block_mem_reg[23][3]  ( .D(n1342), .CLK(clk), .Q(core_block[259])
         );
  DFFPOSX1 \block_mem_reg[23][2]  ( .D(n1341), .CLK(clk), .Q(core_block[258])
         );
  DFFPOSX1 \block_mem_reg[23][1]  ( .D(n1340), .CLK(clk), .Q(core_block[257])
         );
  DFFPOSX1 \block_mem_reg[23][0]  ( .D(n1339), .CLK(clk), .Q(core_block[256])
         );
  DFFPOSX1 \block_mem_reg[24][31]  ( .D(n1338), .CLK(clk), .Q(core_block[255])
         );
  DFFPOSX1 \block_mem_reg[24][30]  ( .D(n1337), .CLK(clk), .Q(core_block[254])
         );
  DFFPOSX1 \block_mem_reg[24][29]  ( .D(n1336), .CLK(clk), .Q(core_block[253])
         );
  DFFPOSX1 \block_mem_reg[24][28]  ( .D(n1335), .CLK(clk), .Q(core_block[252])
         );
  DFFPOSX1 \block_mem_reg[24][27]  ( .D(n1334), .CLK(clk), .Q(core_block[251])
         );
  DFFPOSX1 \block_mem_reg[24][26]  ( .D(n1333), .CLK(clk), .Q(core_block[250])
         );
  DFFPOSX1 \block_mem_reg[24][25]  ( .D(n1332), .CLK(clk), .Q(core_block[249])
         );
  DFFPOSX1 \block_mem_reg[24][24]  ( .D(n1331), .CLK(clk), .Q(core_block[248])
         );
  DFFPOSX1 \block_mem_reg[24][23]  ( .D(n1330), .CLK(clk), .Q(core_block[247])
         );
  DFFPOSX1 \block_mem_reg[24][22]  ( .D(n1329), .CLK(clk), .Q(core_block[246])
         );
  DFFPOSX1 \block_mem_reg[24][21]  ( .D(n1328), .CLK(clk), .Q(core_block[245])
         );
  DFFPOSX1 \block_mem_reg[24][20]  ( .D(n1327), .CLK(clk), .Q(core_block[244])
         );
  DFFPOSX1 \block_mem_reg[24][19]  ( .D(n1326), .CLK(clk), .Q(core_block[243])
         );
  DFFPOSX1 \block_mem_reg[24][18]  ( .D(n1325), .CLK(clk), .Q(core_block[242])
         );
  DFFPOSX1 \block_mem_reg[24][17]  ( .D(n1324), .CLK(clk), .Q(core_block[241])
         );
  DFFPOSX1 \block_mem_reg[24][16]  ( .D(n1323), .CLK(clk), .Q(core_block[240])
         );
  DFFPOSX1 \block_mem_reg[24][15]  ( .D(n1322), .CLK(clk), .Q(core_block[239])
         );
  DFFPOSX1 \block_mem_reg[24][14]  ( .D(n1321), .CLK(clk), .Q(core_block[238])
         );
  DFFPOSX1 \block_mem_reg[24][13]  ( .D(n1320), .CLK(clk), .Q(core_block[237])
         );
  DFFPOSX1 \block_mem_reg[24][12]  ( .D(n1319), .CLK(clk), .Q(core_block[236])
         );
  DFFPOSX1 \block_mem_reg[24][11]  ( .D(n1318), .CLK(clk), .Q(core_block[235])
         );
  DFFPOSX1 \block_mem_reg[24][10]  ( .D(n1317), .CLK(clk), .Q(core_block[234])
         );
  DFFPOSX1 \block_mem_reg[24][9]  ( .D(n1316), .CLK(clk), .Q(core_block[233])
         );
  DFFPOSX1 \block_mem_reg[24][8]  ( .D(n1315), .CLK(clk), .Q(core_block[232])
         );
  DFFPOSX1 \block_mem_reg[24][7]  ( .D(n1314), .CLK(clk), .Q(core_block[231])
         );
  DFFPOSX1 \block_mem_reg[24][6]  ( .D(n1313), .CLK(clk), .Q(core_block[230])
         );
  DFFPOSX1 \block_mem_reg[24][5]  ( .D(n1312), .CLK(clk), .Q(core_block[229])
         );
  DFFPOSX1 \block_mem_reg[24][4]  ( .D(n1311), .CLK(clk), .Q(core_block[228])
         );
  DFFPOSX1 \block_mem_reg[24][3]  ( .D(n1310), .CLK(clk), .Q(core_block[227])
         );
  DFFPOSX1 \block_mem_reg[24][2]  ( .D(n1309), .CLK(clk), .Q(core_block[226])
         );
  DFFPOSX1 \block_mem_reg[24][1]  ( .D(n1308), .CLK(clk), .Q(core_block[225])
         );
  DFFPOSX1 \block_mem_reg[24][0]  ( .D(n1307), .CLK(clk), .Q(core_block[224])
         );
  DFFPOSX1 \block_mem_reg[25][31]  ( .D(n1306), .CLK(clk), .Q(core_block[223])
         );
  DFFPOSX1 \block_mem_reg[25][30]  ( .D(n1305), .CLK(clk), .Q(core_block[222])
         );
  DFFPOSX1 \block_mem_reg[25][29]  ( .D(n1304), .CLK(clk), .Q(core_block[221])
         );
  DFFPOSX1 \block_mem_reg[25][28]  ( .D(n1303), .CLK(clk), .Q(core_block[220])
         );
  DFFPOSX1 \block_mem_reg[25][27]  ( .D(n1302), .CLK(clk), .Q(core_block[219])
         );
  DFFPOSX1 \block_mem_reg[25][26]  ( .D(n1301), .CLK(clk), .Q(core_block[218])
         );
  DFFPOSX1 \block_mem_reg[25][25]  ( .D(n1300), .CLK(clk), .Q(core_block[217])
         );
  DFFPOSX1 \block_mem_reg[25][24]  ( .D(n1299), .CLK(clk), .Q(core_block[216])
         );
  DFFPOSX1 \block_mem_reg[25][23]  ( .D(n1298), .CLK(clk), .Q(core_block[215])
         );
  DFFPOSX1 \block_mem_reg[25][22]  ( .D(n1297), .CLK(clk), .Q(core_block[214])
         );
  DFFPOSX1 \block_mem_reg[25][21]  ( .D(n1296), .CLK(clk), .Q(core_block[213])
         );
  DFFPOSX1 \block_mem_reg[25][20]  ( .D(n1295), .CLK(clk), .Q(core_block[212])
         );
  DFFPOSX1 \block_mem_reg[25][19]  ( .D(n1294), .CLK(clk), .Q(core_block[211])
         );
  DFFPOSX1 \block_mem_reg[25][18]  ( .D(n1293), .CLK(clk), .Q(core_block[210])
         );
  DFFPOSX1 \block_mem_reg[25][17]  ( .D(n1292), .CLK(clk), .Q(core_block[209])
         );
  DFFPOSX1 \block_mem_reg[25][16]  ( .D(n1291), .CLK(clk), .Q(core_block[208])
         );
  DFFPOSX1 \block_mem_reg[25][15]  ( .D(n1290), .CLK(clk), .Q(core_block[207])
         );
  DFFPOSX1 \block_mem_reg[25][14]  ( .D(n1289), .CLK(clk), .Q(core_block[206])
         );
  DFFPOSX1 \block_mem_reg[25][13]  ( .D(n1288), .CLK(clk), .Q(core_block[205])
         );
  DFFPOSX1 \block_mem_reg[25][12]  ( .D(n1287), .CLK(clk), .Q(core_block[204])
         );
  DFFPOSX1 \block_mem_reg[25][11]  ( .D(n1286), .CLK(clk), .Q(core_block[203])
         );
  DFFPOSX1 \block_mem_reg[25][10]  ( .D(n1285), .CLK(clk), .Q(core_block[202])
         );
  DFFPOSX1 \block_mem_reg[25][9]  ( .D(n1284), .CLK(clk), .Q(core_block[201])
         );
  DFFPOSX1 \block_mem_reg[25][8]  ( .D(n1283), .CLK(clk), .Q(core_block[200])
         );
  DFFPOSX1 \block_mem_reg[25][7]  ( .D(n1282), .CLK(clk), .Q(core_block[199])
         );
  DFFPOSX1 \block_mem_reg[25][6]  ( .D(n1281), .CLK(clk), .Q(core_block[198])
         );
  DFFPOSX1 \block_mem_reg[25][5]  ( .D(n1280), .CLK(clk), .Q(core_block[197])
         );
  DFFPOSX1 \block_mem_reg[25][4]  ( .D(n1279), .CLK(clk), .Q(core_block[196])
         );
  DFFPOSX1 \block_mem_reg[25][3]  ( .D(n1278), .CLK(clk), .Q(core_block[195])
         );
  DFFPOSX1 \block_mem_reg[25][2]  ( .D(n1277), .CLK(clk), .Q(core_block[194])
         );
  DFFPOSX1 \block_mem_reg[25][1]  ( .D(n1276), .CLK(clk), .Q(core_block[193])
         );
  DFFPOSX1 \block_mem_reg[25][0]  ( .D(n1275), .CLK(clk), .Q(core_block[192])
         );
  DFFPOSX1 \block_mem_reg[26][31]  ( .D(n1274), .CLK(clk), .Q(core_block[191])
         );
  DFFPOSX1 \block_mem_reg[26][30]  ( .D(n1273), .CLK(clk), .Q(core_block[190])
         );
  DFFPOSX1 \block_mem_reg[26][29]  ( .D(n1272), .CLK(clk), .Q(core_block[189])
         );
  DFFPOSX1 \block_mem_reg[26][28]  ( .D(n1271), .CLK(clk), .Q(core_block[188])
         );
  DFFPOSX1 \block_mem_reg[26][27]  ( .D(n1270), .CLK(clk), .Q(core_block[187])
         );
  DFFPOSX1 \block_mem_reg[26][26]  ( .D(n1269), .CLK(clk), .Q(core_block[186])
         );
  DFFPOSX1 \block_mem_reg[26][25]  ( .D(n1268), .CLK(clk), .Q(core_block[185])
         );
  DFFPOSX1 \block_mem_reg[26][24]  ( .D(n1267), .CLK(clk), .Q(core_block[184])
         );
  DFFPOSX1 \block_mem_reg[26][23]  ( .D(n1266), .CLK(clk), .Q(core_block[183])
         );
  DFFPOSX1 \block_mem_reg[26][22]  ( .D(n1265), .CLK(clk), .Q(core_block[182])
         );
  DFFPOSX1 \block_mem_reg[26][21]  ( .D(n1264), .CLK(clk), .Q(core_block[181])
         );
  DFFPOSX1 \block_mem_reg[26][20]  ( .D(n1263), .CLK(clk), .Q(core_block[180])
         );
  DFFPOSX1 \block_mem_reg[26][19]  ( .D(n1262), .CLK(clk), .Q(core_block[179])
         );
  DFFPOSX1 \block_mem_reg[26][18]  ( .D(n1261), .CLK(clk), .Q(core_block[178])
         );
  DFFPOSX1 \block_mem_reg[26][17]  ( .D(n1260), .CLK(clk), .Q(core_block[177])
         );
  DFFPOSX1 \block_mem_reg[26][16]  ( .D(n1259), .CLK(clk), .Q(core_block[176])
         );
  DFFPOSX1 \block_mem_reg[26][15]  ( .D(n1258), .CLK(clk), .Q(core_block[175])
         );
  DFFPOSX1 \block_mem_reg[26][14]  ( .D(n1257), .CLK(clk), .Q(core_block[174])
         );
  DFFPOSX1 \block_mem_reg[26][13]  ( .D(n1256), .CLK(clk), .Q(core_block[173])
         );
  DFFPOSX1 \block_mem_reg[26][12]  ( .D(n1255), .CLK(clk), .Q(core_block[172])
         );
  DFFPOSX1 \block_mem_reg[26][11]  ( .D(n1254), .CLK(clk), .Q(core_block[171])
         );
  DFFPOSX1 \block_mem_reg[26][10]  ( .D(n1253), .CLK(clk), .Q(core_block[170])
         );
  DFFPOSX1 \block_mem_reg[26][9]  ( .D(n1252), .CLK(clk), .Q(core_block[169])
         );
  DFFPOSX1 \block_mem_reg[26][8]  ( .D(n1251), .CLK(clk), .Q(core_block[168])
         );
  DFFPOSX1 \block_mem_reg[26][7]  ( .D(n1250), .CLK(clk), .Q(core_block[167])
         );
  DFFPOSX1 \block_mem_reg[26][6]  ( .D(n1249), .CLK(clk), .Q(core_block[166])
         );
  DFFPOSX1 \block_mem_reg[26][5]  ( .D(n1248), .CLK(clk), .Q(core_block[165])
         );
  DFFPOSX1 \block_mem_reg[26][4]  ( .D(n1247), .CLK(clk), .Q(core_block[164])
         );
  DFFPOSX1 \block_mem_reg[26][3]  ( .D(n1246), .CLK(clk), .Q(core_block[163])
         );
  DFFPOSX1 \block_mem_reg[26][2]  ( .D(n1245), .CLK(clk), .Q(core_block[162])
         );
  DFFPOSX1 \block_mem_reg[26][1]  ( .D(n1244), .CLK(clk), .Q(core_block[161])
         );
  DFFPOSX1 \block_mem_reg[26][0]  ( .D(n1243), .CLK(clk), .Q(core_block[160])
         );
  DFFPOSX1 \block_mem_reg[27][31]  ( .D(n1242), .CLK(clk), .Q(core_block[159])
         );
  DFFPOSX1 \block_mem_reg[27][30]  ( .D(n1241), .CLK(clk), .Q(core_block[158])
         );
  DFFPOSX1 \block_mem_reg[27][29]  ( .D(n1240), .CLK(clk), .Q(core_block[157])
         );
  DFFPOSX1 \block_mem_reg[27][28]  ( .D(n1239), .CLK(clk), .Q(core_block[156])
         );
  DFFPOSX1 \block_mem_reg[27][27]  ( .D(n1238), .CLK(clk), .Q(core_block[155])
         );
  DFFPOSX1 \block_mem_reg[27][26]  ( .D(n1237), .CLK(clk), .Q(core_block[154])
         );
  DFFPOSX1 \block_mem_reg[27][25]  ( .D(n1236), .CLK(clk), .Q(core_block[153])
         );
  DFFPOSX1 \block_mem_reg[27][24]  ( .D(n1235), .CLK(clk), .Q(core_block[152])
         );
  DFFPOSX1 \block_mem_reg[27][23]  ( .D(n1234), .CLK(clk), .Q(core_block[151])
         );
  DFFPOSX1 \block_mem_reg[27][22]  ( .D(n1233), .CLK(clk), .Q(core_block[150])
         );
  DFFPOSX1 \block_mem_reg[27][21]  ( .D(n1232), .CLK(clk), .Q(core_block[149])
         );
  DFFPOSX1 \block_mem_reg[27][20]  ( .D(n1231), .CLK(clk), .Q(core_block[148])
         );
  DFFPOSX1 \block_mem_reg[27][19]  ( .D(n1230), .CLK(clk), .Q(core_block[147])
         );
  DFFPOSX1 \block_mem_reg[27][18]  ( .D(n1229), .CLK(clk), .Q(core_block[146])
         );
  DFFPOSX1 \block_mem_reg[27][17]  ( .D(n1228), .CLK(clk), .Q(core_block[145])
         );
  DFFPOSX1 \block_mem_reg[27][16]  ( .D(n1227), .CLK(clk), .Q(core_block[144])
         );
  DFFPOSX1 \block_mem_reg[27][15]  ( .D(n1226), .CLK(clk), .Q(core_block[143])
         );
  DFFPOSX1 \block_mem_reg[27][14]  ( .D(n1225), .CLK(clk), .Q(core_block[142])
         );
  DFFPOSX1 \block_mem_reg[27][13]  ( .D(n1224), .CLK(clk), .Q(core_block[141])
         );
  DFFPOSX1 \block_mem_reg[27][12]  ( .D(n1223), .CLK(clk), .Q(core_block[140])
         );
  DFFPOSX1 \block_mem_reg[27][11]  ( .D(n1222), .CLK(clk), .Q(core_block[139])
         );
  DFFPOSX1 \block_mem_reg[27][10]  ( .D(n1221), .CLK(clk), .Q(core_block[138])
         );
  DFFPOSX1 \block_mem_reg[27][9]  ( .D(n1220), .CLK(clk), .Q(core_block[137])
         );
  DFFPOSX1 \block_mem_reg[27][8]  ( .D(n1219), .CLK(clk), .Q(core_block[136])
         );
  DFFPOSX1 \block_mem_reg[27][7]  ( .D(n1218), .CLK(clk), .Q(core_block[135])
         );
  DFFPOSX1 \block_mem_reg[27][6]  ( .D(n1217), .CLK(clk), .Q(core_block[134])
         );
  DFFPOSX1 \block_mem_reg[27][5]  ( .D(n1216), .CLK(clk), .Q(core_block[133])
         );
  DFFPOSX1 \block_mem_reg[27][4]  ( .D(n1215), .CLK(clk), .Q(core_block[132])
         );
  DFFPOSX1 \block_mem_reg[27][3]  ( .D(n1214), .CLK(clk), .Q(core_block[131])
         );
  DFFPOSX1 \block_mem_reg[27][2]  ( .D(n1213), .CLK(clk), .Q(core_block[130])
         );
  DFFPOSX1 \block_mem_reg[27][1]  ( .D(n1212), .CLK(clk), .Q(core_block[129])
         );
  DFFPOSX1 \block_mem_reg[27][0]  ( .D(n1211), .CLK(clk), .Q(core_block[128])
         );
  DFFPOSX1 \block_mem_reg[28][31]  ( .D(n1210), .CLK(clk), .Q(core_block[127])
         );
  DFFPOSX1 \block_mem_reg[28][30]  ( .D(n1209), .CLK(clk), .Q(core_block[126])
         );
  DFFPOSX1 \block_mem_reg[28][29]  ( .D(n1208), .CLK(clk), .Q(core_block[125])
         );
  DFFPOSX1 \block_mem_reg[28][28]  ( .D(n1207), .CLK(clk), .Q(core_block[124])
         );
  DFFPOSX1 \block_mem_reg[28][27]  ( .D(n1206), .CLK(clk), .Q(core_block[123])
         );
  DFFPOSX1 \block_mem_reg[28][26]  ( .D(n1205), .CLK(clk), .Q(core_block[122])
         );
  DFFPOSX1 \block_mem_reg[28][25]  ( .D(n1204), .CLK(clk), .Q(core_block[121])
         );
  DFFPOSX1 \block_mem_reg[28][24]  ( .D(n1203), .CLK(clk), .Q(core_block[120])
         );
  DFFPOSX1 \block_mem_reg[28][23]  ( .D(n1202), .CLK(clk), .Q(core_block[119])
         );
  DFFPOSX1 \block_mem_reg[28][22]  ( .D(n1201), .CLK(clk), .Q(core_block[118])
         );
  DFFPOSX1 \block_mem_reg[28][21]  ( .D(n1200), .CLK(clk), .Q(core_block[117])
         );
  DFFPOSX1 \block_mem_reg[28][20]  ( .D(n1199), .CLK(clk), .Q(core_block[116])
         );
  DFFPOSX1 \block_mem_reg[28][19]  ( .D(n1198), .CLK(clk), .Q(core_block[115])
         );
  DFFPOSX1 \block_mem_reg[28][18]  ( .D(n1197), .CLK(clk), .Q(core_block[114])
         );
  DFFPOSX1 \block_mem_reg[28][17]  ( .D(n1196), .CLK(clk), .Q(core_block[113])
         );
  DFFPOSX1 \block_mem_reg[28][16]  ( .D(n1195), .CLK(clk), .Q(core_block[112])
         );
  DFFPOSX1 \block_mem_reg[28][15]  ( .D(n1194), .CLK(clk), .Q(core_block[111])
         );
  DFFPOSX1 \block_mem_reg[28][14]  ( .D(n1193), .CLK(clk), .Q(core_block[110])
         );
  DFFPOSX1 \block_mem_reg[28][13]  ( .D(n1192), .CLK(clk), .Q(core_block[109])
         );
  DFFPOSX1 \block_mem_reg[28][12]  ( .D(n1191), .CLK(clk), .Q(core_block[108])
         );
  DFFPOSX1 \block_mem_reg[28][11]  ( .D(n1190), .CLK(clk), .Q(core_block[107])
         );
  DFFPOSX1 \block_mem_reg[28][10]  ( .D(n1189), .CLK(clk), .Q(core_block[106])
         );
  DFFPOSX1 \block_mem_reg[28][9]  ( .D(n1188), .CLK(clk), .Q(core_block[105])
         );
  DFFPOSX1 \block_mem_reg[28][8]  ( .D(n1187), .CLK(clk), .Q(core_block[104])
         );
  DFFPOSX1 \block_mem_reg[28][7]  ( .D(n1186), .CLK(clk), .Q(core_block[103])
         );
  DFFPOSX1 \block_mem_reg[28][6]  ( .D(n1185), .CLK(clk), .Q(core_block[102])
         );
  DFFPOSX1 \block_mem_reg[28][5]  ( .D(n1184), .CLK(clk), .Q(core_block[101])
         );
  DFFPOSX1 \block_mem_reg[28][4]  ( .D(n1183), .CLK(clk), .Q(core_block[100])
         );
  DFFPOSX1 \block_mem_reg[28][3]  ( .D(n1182), .CLK(clk), .Q(core_block[99])
         );
  DFFPOSX1 \block_mem_reg[28][2]  ( .D(n1181), .CLK(clk), .Q(core_block[98])
         );
  DFFPOSX1 \block_mem_reg[28][1]  ( .D(n1180), .CLK(clk), .Q(core_block[97])
         );
  DFFPOSX1 \block_mem_reg[28][0]  ( .D(n1179), .CLK(clk), .Q(core_block[96])
         );
  DFFPOSX1 \block_mem_reg[29][31]  ( .D(n1178), .CLK(clk), .Q(core_block[95])
         );
  DFFPOSX1 \block_mem_reg[29][30]  ( .D(n1177), .CLK(clk), .Q(core_block[94])
         );
  DFFPOSX1 \block_mem_reg[29][29]  ( .D(n1176), .CLK(clk), .Q(core_block[93])
         );
  DFFPOSX1 \block_mem_reg[29][28]  ( .D(n1175), .CLK(clk), .Q(core_block[92])
         );
  DFFPOSX1 \block_mem_reg[29][27]  ( .D(n1174), .CLK(clk), .Q(core_block[91])
         );
  DFFPOSX1 \block_mem_reg[29][26]  ( .D(n1173), .CLK(clk), .Q(core_block[90])
         );
  DFFPOSX1 \block_mem_reg[29][25]  ( .D(n1172), .CLK(clk), .Q(core_block[89])
         );
  DFFPOSX1 \block_mem_reg[29][24]  ( .D(n1171), .CLK(clk), .Q(core_block[88])
         );
  DFFPOSX1 \block_mem_reg[29][23]  ( .D(n1170), .CLK(clk), .Q(core_block[87])
         );
  DFFPOSX1 \block_mem_reg[29][22]  ( .D(n1169), .CLK(clk), .Q(core_block[86])
         );
  DFFPOSX1 \block_mem_reg[29][21]  ( .D(n1168), .CLK(clk), .Q(core_block[85])
         );
  DFFPOSX1 \block_mem_reg[29][20]  ( .D(n1167), .CLK(clk), .Q(core_block[84])
         );
  DFFPOSX1 \block_mem_reg[29][19]  ( .D(n1166), .CLK(clk), .Q(core_block[83])
         );
  DFFPOSX1 \block_mem_reg[29][18]  ( .D(n1165), .CLK(clk), .Q(core_block[82])
         );
  DFFPOSX1 \block_mem_reg[29][17]  ( .D(n1164), .CLK(clk), .Q(core_block[81])
         );
  DFFPOSX1 \block_mem_reg[29][16]  ( .D(n1163), .CLK(clk), .Q(core_block[80])
         );
  DFFPOSX1 \block_mem_reg[29][15]  ( .D(n1162), .CLK(clk), .Q(core_block[79])
         );
  DFFPOSX1 \block_mem_reg[29][14]  ( .D(n1161), .CLK(clk), .Q(core_block[78])
         );
  DFFPOSX1 \block_mem_reg[29][13]  ( .D(n1160), .CLK(clk), .Q(core_block[77])
         );
  DFFPOSX1 \block_mem_reg[29][12]  ( .D(n1159), .CLK(clk), .Q(core_block[76])
         );
  DFFPOSX1 \block_mem_reg[29][11]  ( .D(n1158), .CLK(clk), .Q(core_block[75])
         );
  DFFPOSX1 \block_mem_reg[29][10]  ( .D(n1157), .CLK(clk), .Q(core_block[74])
         );
  DFFPOSX1 \block_mem_reg[29][9]  ( .D(n1156), .CLK(clk), .Q(core_block[73])
         );
  DFFPOSX1 \block_mem_reg[29][8]  ( .D(n1155), .CLK(clk), .Q(core_block[72])
         );
  DFFPOSX1 \block_mem_reg[29][7]  ( .D(n1154), .CLK(clk), .Q(core_block[71])
         );
  DFFPOSX1 \block_mem_reg[29][6]  ( .D(n1153), .CLK(clk), .Q(core_block[70])
         );
  DFFPOSX1 \block_mem_reg[29][5]  ( .D(n1152), .CLK(clk), .Q(core_block[69])
         );
  DFFPOSX1 \block_mem_reg[29][4]  ( .D(n1151), .CLK(clk), .Q(core_block[68])
         );
  DFFPOSX1 \block_mem_reg[29][3]  ( .D(n1150), .CLK(clk), .Q(core_block[67])
         );
  DFFPOSX1 \block_mem_reg[29][2]  ( .D(n1149), .CLK(clk), .Q(core_block[66])
         );
  DFFPOSX1 \block_mem_reg[29][1]  ( .D(n1148), .CLK(clk), .Q(core_block[65])
         );
  DFFPOSX1 \block_mem_reg[29][0]  ( .D(n1147), .CLK(clk), .Q(core_block[64])
         );
  DFFPOSX1 \block_mem_reg[30][31]  ( .D(n1146), .CLK(clk), .Q(core_block[63])
         );
  DFFPOSX1 \block_mem_reg[30][30]  ( .D(n1145), .CLK(clk), .Q(core_block[62])
         );
  DFFPOSX1 \block_mem_reg[30][29]  ( .D(n1144), .CLK(clk), .Q(core_block[61])
         );
  DFFPOSX1 \block_mem_reg[30][28]  ( .D(n1143), .CLK(clk), .Q(core_block[60])
         );
  DFFPOSX1 \block_mem_reg[30][27]  ( .D(n1142), .CLK(clk), .Q(core_block[59])
         );
  DFFPOSX1 \block_mem_reg[30][26]  ( .D(n1141), .CLK(clk), .Q(core_block[58])
         );
  DFFPOSX1 \block_mem_reg[30][25]  ( .D(n1140), .CLK(clk), .Q(core_block[57])
         );
  DFFPOSX1 \block_mem_reg[30][24]  ( .D(n1139), .CLK(clk), .Q(core_block[56])
         );
  DFFPOSX1 \block_mem_reg[30][23]  ( .D(n1138), .CLK(clk), .Q(core_block[55])
         );
  DFFPOSX1 \block_mem_reg[30][22]  ( .D(n1137), .CLK(clk), .Q(core_block[54])
         );
  DFFPOSX1 \block_mem_reg[30][21]  ( .D(n1136), .CLK(clk), .Q(core_block[53])
         );
  DFFPOSX1 \block_mem_reg[30][20]  ( .D(n1135), .CLK(clk), .Q(core_block[52])
         );
  DFFPOSX1 \block_mem_reg[30][19]  ( .D(n1134), .CLK(clk), .Q(core_block[51])
         );
  DFFPOSX1 \block_mem_reg[30][18]  ( .D(n1133), .CLK(clk), .Q(core_block[50])
         );
  DFFPOSX1 \block_mem_reg[30][17]  ( .D(n1132), .CLK(clk), .Q(core_block[49])
         );
  DFFPOSX1 \block_mem_reg[30][16]  ( .D(n1131), .CLK(clk), .Q(core_block[48])
         );
  DFFPOSX1 \block_mem_reg[30][15]  ( .D(n1130), .CLK(clk), .Q(core_block[47])
         );
  DFFPOSX1 \block_mem_reg[30][14]  ( .D(n1129), .CLK(clk), .Q(core_block[46])
         );
  DFFPOSX1 \block_mem_reg[30][13]  ( .D(n1128), .CLK(clk), .Q(core_block[45])
         );
  DFFPOSX1 \block_mem_reg[30][12]  ( .D(n1127), .CLK(clk), .Q(core_block[44])
         );
  DFFPOSX1 \block_mem_reg[30][11]  ( .D(n1126), .CLK(clk), .Q(core_block[43])
         );
  DFFPOSX1 \block_mem_reg[30][10]  ( .D(n1125), .CLK(clk), .Q(core_block[42])
         );
  DFFPOSX1 \block_mem_reg[30][9]  ( .D(n1124), .CLK(clk), .Q(core_block[41])
         );
  DFFPOSX1 \block_mem_reg[30][8]  ( .D(n1123), .CLK(clk), .Q(core_block[40])
         );
  DFFPOSX1 \block_mem_reg[30][7]  ( .D(n1122), .CLK(clk), .Q(core_block[39])
         );
  DFFPOSX1 \block_mem_reg[30][6]  ( .D(n1121), .CLK(clk), .Q(core_block[38])
         );
  DFFPOSX1 \block_mem_reg[30][5]  ( .D(n1120), .CLK(clk), .Q(core_block[37])
         );
  DFFPOSX1 \block_mem_reg[30][4]  ( .D(n1119), .CLK(clk), .Q(core_block[36])
         );
  DFFPOSX1 \block_mem_reg[30][3]  ( .D(n1118), .CLK(clk), .Q(core_block[35])
         );
  DFFPOSX1 \block_mem_reg[30][2]  ( .D(n1117), .CLK(clk), .Q(core_block[34])
         );
  DFFPOSX1 \block_mem_reg[30][1]  ( .D(n1116), .CLK(clk), .Q(core_block[33])
         );
  DFFPOSX1 \block_mem_reg[30][0]  ( .D(n1115), .CLK(clk), .Q(core_block[32])
         );
  DFFPOSX1 \block_mem_reg[31][31]  ( .D(n1114), .CLK(clk), .Q(core_block[31])
         );
  DFFPOSX1 \block_mem_reg[31][30]  ( .D(n1113), .CLK(clk), .Q(core_block[30])
         );
  DFFPOSX1 \block_mem_reg[31][29]  ( .D(n1112), .CLK(clk), .Q(core_block[29])
         );
  DFFPOSX1 \block_mem_reg[31][28]  ( .D(n1111), .CLK(clk), .Q(core_block[28])
         );
  DFFPOSX1 \block_mem_reg[31][27]  ( .D(n1110), .CLK(clk), .Q(core_block[27])
         );
  DFFPOSX1 \block_mem_reg[31][26]  ( .D(n1109), .CLK(clk), .Q(core_block[26])
         );
  DFFPOSX1 \block_mem_reg[31][25]  ( .D(n1108), .CLK(clk), .Q(core_block[25])
         );
  DFFPOSX1 \block_mem_reg[31][24]  ( .D(n1107), .CLK(clk), .Q(core_block[24])
         );
  DFFPOSX1 \block_mem_reg[31][23]  ( .D(n1106), .CLK(clk), .Q(core_block[23])
         );
  DFFPOSX1 \block_mem_reg[31][22]  ( .D(n1105), .CLK(clk), .Q(core_block[22])
         );
  DFFPOSX1 \block_mem_reg[31][21]  ( .D(n1104), .CLK(clk), .Q(core_block[21])
         );
  DFFPOSX1 \block_mem_reg[31][20]  ( .D(n1103), .CLK(clk), .Q(core_block[20])
         );
  DFFPOSX1 \block_mem_reg[31][19]  ( .D(n1102), .CLK(clk), .Q(core_block[19])
         );
  DFFPOSX1 \block_mem_reg[31][18]  ( .D(n1101), .CLK(clk), .Q(core_block[18])
         );
  DFFPOSX1 \block_mem_reg[31][17]  ( .D(n1100), .CLK(clk), .Q(core_block[17])
         );
  DFFPOSX1 \block_mem_reg[31][16]  ( .D(n1099), .CLK(clk), .Q(core_block[16])
         );
  DFFPOSX1 \block_mem_reg[31][15]  ( .D(n1098), .CLK(clk), .Q(core_block[15])
         );
  DFFPOSX1 \block_mem_reg[31][14]  ( .D(n1097), .CLK(clk), .Q(core_block[14])
         );
  DFFPOSX1 \block_mem_reg[31][13]  ( .D(n1096), .CLK(clk), .Q(core_block[13])
         );
  DFFPOSX1 \block_mem_reg[31][12]  ( .D(n1095), .CLK(clk), .Q(core_block[12])
         );
  DFFPOSX1 \block_mem_reg[31][11]  ( .D(n1094), .CLK(clk), .Q(core_block[11])
         );
  DFFPOSX1 \block_mem_reg[31][10]  ( .D(n1093), .CLK(clk), .Q(core_block[10])
         );
  DFFPOSX1 \block_mem_reg[31][9]  ( .D(n1092), .CLK(clk), .Q(core_block[9]) );
  DFFPOSX1 \block_mem_reg[31][8]  ( .D(n1091), .CLK(clk), .Q(core_block[8]) );
  DFFPOSX1 \block_mem_reg[31][7]  ( .D(n1090), .CLK(clk), .Q(core_block[7]) );
  DFFPOSX1 \block_mem_reg[31][6]  ( .D(n1089), .CLK(clk), .Q(core_block[6]) );
  DFFPOSX1 \block_mem_reg[31][5]  ( .D(n1088), .CLK(clk), .Q(core_block[5]) );
  DFFPOSX1 \block_mem_reg[31][4]  ( .D(n1087), .CLK(clk), .Q(core_block[4]) );
  DFFPOSX1 \block_mem_reg[31][3]  ( .D(n1086), .CLK(clk), .Q(core_block[3]) );
  DFFPOSX1 \block_mem_reg[31][2]  ( .D(n1085), .CLK(clk), .Q(core_block[2]) );
  DFFPOSX1 \block_mem_reg[31][1]  ( .D(n1084), .CLK(clk), .Q(core_block[1]) );
  DFFPOSX1 \block_mem_reg[31][0]  ( .D(n1083), .CLK(clk), .Q(core_block[0]) );
  DFFPOSX1 init_reg_reg ( .D(n2170), .CLK(clk), .Q(core_init) );
  DFFPOSX1 digest_valid_reg_reg ( .D(N62), .CLK(clk), .Q(digest_valid_reg) );
  DFFPOSX1 ready_reg_reg ( .D(N61), .CLK(clk), .Q(ready_reg) );
  NAND2X1 U3 ( .A(n5), .B(n6), .Y(read_data_30) );
  OAI21X1 U6 ( .A(n7), .B(n8), .C(n5), .Y(read_data_1) );
  AOI22X1 U7 ( .A(core_next), .B(N159), .C(digest_valid_reg), .D(N162), .Y(n7)
         );
  OAI21X1 U8 ( .A(n9), .B(n8), .C(n5), .Y(read_data_0) );
  INVX1 U9 ( .A(read_data_6), .Y(n5) );
  AOI22X1 U10 ( .A(core_init), .B(N159), .C(ready_reg), .D(N162), .Y(n9) );
  NOR2X1 U11 ( .A(n10), .B(n11), .Y(read_data_6) );
  INVX1 U12 ( .A(n12), .Y(read_data_5) );
  OAI21X1 U13 ( .A(n13), .B(n14), .C(cs), .Y(n12) );
  AND2X1 U14 ( .A(n15), .B(N152), .Y(n13) );
  AND2X1 U15 ( .A(cs), .B(n14), .Y(read_data_8) );
  OAI21X1 U16 ( .A(n16), .B(n17), .C(n10), .Y(n14) );
  NAND3X1 U17 ( .A(n15), .B(n18), .C(N148), .Y(n10) );
  OR2X1 U18 ( .A(read_data_4), .B(read_data_26), .Y(read_data[17]) );
  INVX1 U19 ( .A(n6), .Y(read_data_26) );
  NAND2X1 U20 ( .A(n19), .B(N152), .Y(n6) );
  NOR2X1 U21 ( .A(n8), .B(n17), .Y(read_data_4) );
  INVX1 U22 ( .A(N155), .Y(n17) );
  INVX1 U23 ( .A(n19), .Y(n8) );
  OAI21X1 U24 ( .A(n11), .B(n20), .C(n21), .Y(error) );
  NAND2X1 U25 ( .A(N165), .B(n19), .Y(n21) );
  NOR2X1 U26 ( .A(n11), .B(n16), .Y(n19) );
  INVX1 U27 ( .A(n15), .Y(n16) );
  NOR2X1 U28 ( .A(n22), .B(we), .Y(n15) );
  NAND2X1 U29 ( .A(n22), .B(n23), .Y(n20) );
  INVX1 U30 ( .A(we), .Y(n23) );
  NAND2X1 U31 ( .A(N144), .B(N200), .Y(n22) );
  INVX1 U32 ( .A(cs), .Y(n11) );
  OAI21X1 U33 ( .A(n2168), .B(n25), .C(reset_n), .Y(N99) );
  INVX1 U34 ( .A(N219), .Y(n25) );
  OAI21X1 U35 ( .A(n2168), .B(n26), .C(reset_n), .Y(N98) );
  INVX1 U36 ( .A(N218), .Y(n26) );
  OAI21X1 U37 ( .A(n2168), .B(n27), .C(reset_n), .Y(N97) );
  INVX1 U38 ( .A(N217), .Y(n27) );
  OAI21X1 U39 ( .A(n2168), .B(n28), .C(reset_n), .Y(N96) );
  INVX1 U40 ( .A(N216), .Y(n28) );
  OAI21X1 U41 ( .A(n2168), .B(n29), .C(reset_n), .Y(N95) );
  INVX1 U42 ( .A(N215), .Y(n29) );
  OAI21X1 U43 ( .A(n2168), .B(n30), .C(reset_n), .Y(N94) );
  INVX1 U44 ( .A(N214), .Y(n30) );
  AND2X1 U45 ( .A(write_data[31]), .B(reset_n), .Y(N93) );
  AND2X1 U46 ( .A(write_data[30]), .B(reset_n), .Y(N92) );
  AND2X1 U47 ( .A(write_data[29]), .B(reset_n), .Y(N91) );
  AND2X1 U48 ( .A(write_data[28]), .B(reset_n), .Y(N90) );
  AND2X1 U49 ( .A(write_data[27]), .B(reset_n), .Y(N89) );
  AND2X1 U50 ( .A(write_data[26]), .B(reset_n), .Y(N88) );
  AND2X1 U51 ( .A(write_data[25]), .B(reset_n), .Y(N87) );
  AND2X1 U52 ( .A(write_data[24]), .B(reset_n), .Y(N86) );
  AND2X1 U53 ( .A(write_data[23]), .B(reset_n), .Y(N85) );
  AND2X1 U54 ( .A(write_data[22]), .B(reset_n), .Y(N84) );
  AND2X1 U55 ( .A(write_data[21]), .B(reset_n), .Y(N83) );
  AND2X1 U56 ( .A(write_data[20]), .B(reset_n), .Y(N82) );
  AND2X1 U57 ( .A(write_data[19]), .B(reset_n), .Y(N81) );
  AND2X1 U58 ( .A(write_data[18]), .B(reset_n), .Y(N80) );
  AND2X1 U59 ( .A(write_data[17]), .B(reset_n), .Y(N79) );
  AND2X1 U60 ( .A(write_data[16]), .B(reset_n), .Y(N78) );
  AND2X1 U61 ( .A(write_data[15]), .B(reset_n), .Y(N77) );
  AND2X1 U62 ( .A(write_data[14]), .B(reset_n), .Y(N76) );
  AND2X1 U63 ( .A(write_data[13]), .B(reset_n), .Y(N75) );
  AND2X1 U64 ( .A(write_data[12]), .B(reset_n), .Y(N74) );
  AND2X1 U65 ( .A(write_data[11]), .B(reset_n), .Y(N73) );
  AND2X1 U66 ( .A(write_data[10]), .B(reset_n), .Y(N72) );
  AND2X1 U67 ( .A(write_data[9]), .B(reset_n), .Y(N71) );
  AND2X1 U68 ( .A(write_data[8]), .B(reset_n), .Y(N70) );
  AND2X1 U69 ( .A(write_data[7]), .B(reset_n), .Y(N69) );
  AND2X1 U70 ( .A(write_data[6]), .B(reset_n), .Y(N68) );
  AND2X1 U71 ( .A(write_data[5]), .B(reset_n), .Y(N67) );
  AND2X1 U72 ( .A(write_data[4]), .B(reset_n), .Y(N66) );
  AND2X1 U73 ( .A(write_data[3]), .B(reset_n), .Y(N65) );
  AND2X1 U74 ( .A(write_data[2]), .B(reset_n), .Y(N64) );
  OAI21X1 U75 ( .A(n2168), .B(n31), .C(reset_n), .Y(N63) );
  INVX1 U76 ( .A(N213), .Y(n31) );
  AND2X1 U77 ( .A(core_digest_valid), .B(reset_n), .Y(N62) );
  AND2X1 U78 ( .A(core_ready), .B(reset_n), .Y(N61) );
  AND2X1 U79 ( .A(write_data[1]), .B(reset_n), .Y(N60) );
  AND2X1 U80 ( .A(write_data[0]), .B(reset_n), .Y(N59) );
  NOR2X1 U81 ( .A(n32), .B(N0), .Y(N164) );
  NOR2X1 U82 ( .A(n32), .B(n18), .Y(N163) );
  INVX1 U83 ( .A(address[1]), .Y(n32) );
  NAND2X1 U84 ( .A(address[0]), .B(n33), .Y(N161) );
  NAND2X1 U85 ( .A(n18), .B(n33), .Y(N158) );
  INVX1 U86 ( .A(N157), .Y(n33) );
  OR2X1 U87 ( .A(N153), .B(address[0]), .Y(N154) );
  OR2X1 U88 ( .A(N150), .B(n18), .Y(N151) );
  INVX1 U89 ( .A(address[0]), .Y(n18) );
  OAI21X1 U90 ( .A(n2168), .B(n34), .C(reset_n), .Y(N124) );
  INVX1 U91 ( .A(N244), .Y(n34) );
  OAI21X1 U92 ( .A(n2168), .B(n35), .C(reset_n), .Y(N123) );
  INVX1 U93 ( .A(N243), .Y(n35) );
  OAI21X1 U94 ( .A(n2168), .B(n36), .C(reset_n), .Y(N122) );
  INVX1 U95 ( .A(N242), .Y(n36) );
  OAI21X1 U96 ( .A(n2168), .B(n37), .C(reset_n), .Y(N121) );
  INVX1 U97 ( .A(N241), .Y(n37) );
  OAI21X1 U98 ( .A(n2168), .B(n38), .C(reset_n), .Y(N120) );
  INVX1 U99 ( .A(N240), .Y(n38) );
  OAI21X1 U100 ( .A(n2168), .B(n39), .C(reset_n), .Y(N119) );
  INVX1 U101 ( .A(N239), .Y(n39) );
  OAI21X1 U102 ( .A(n2168), .B(n40), .C(reset_n), .Y(N118) );
  INVX1 U103 ( .A(N238), .Y(n40) );
  OAI21X1 U104 ( .A(n2168), .B(n41), .C(reset_n), .Y(N117) );
  INVX1 U105 ( .A(N237), .Y(n41) );
  OAI21X1 U106 ( .A(n2168), .B(n42), .C(reset_n), .Y(N116) );
  INVX1 U107 ( .A(N236), .Y(n42) );
  OAI21X1 U108 ( .A(n2168), .B(n43), .C(reset_n), .Y(N115) );
  INVX1 U109 ( .A(N235), .Y(n43) );
  OAI21X1 U110 ( .A(n2168), .B(n44), .C(reset_n), .Y(N114) );
  INVX1 U111 ( .A(N234), .Y(n44) );
  OAI21X1 U112 ( .A(n2168), .B(n45), .C(reset_n), .Y(N113) );
  INVX1 U113 ( .A(N233), .Y(n45) );
  OAI21X1 U114 ( .A(n2168), .B(n46), .C(reset_n), .Y(N112) );
  INVX1 U115 ( .A(N232), .Y(n46) );
  OAI21X1 U116 ( .A(n2168), .B(n47), .C(reset_n), .Y(N111) );
  INVX1 U117 ( .A(N231), .Y(n47) );
  OAI21X1 U118 ( .A(n2168), .B(n48), .C(reset_n), .Y(N110) );
  INVX1 U119 ( .A(N230), .Y(n48) );
  OAI21X1 U120 ( .A(n2168), .B(n49), .C(reset_n), .Y(N109) );
  INVX1 U121 ( .A(N229), .Y(n49) );
  OAI21X1 U122 ( .A(n2168), .B(n50), .C(reset_n), .Y(N108) );
  INVX1 U123 ( .A(N228), .Y(n50) );
  OAI21X1 U124 ( .A(n2168), .B(n51), .C(reset_n), .Y(N107) );
  INVX1 U125 ( .A(N227), .Y(n51) );
  OAI21X1 U126 ( .A(n2168), .B(n52), .C(reset_n), .Y(N106) );
  INVX1 U127 ( .A(N226), .Y(n52) );
  OAI21X1 U128 ( .A(n2168), .B(n53), .C(reset_n), .Y(N105) );
  INVX1 U129 ( .A(N225), .Y(n53) );
  OAI21X1 U130 ( .A(n2168), .B(n54), .C(reset_n), .Y(N104) );
  INVX1 U131 ( .A(N224), .Y(n54) );
  OAI21X1 U132 ( .A(n2168), .B(n55), .C(reset_n), .Y(N103) );
  INVX1 U133 ( .A(N223), .Y(n55) );
  OAI21X1 U134 ( .A(n2168), .B(n56), .C(reset_n), .Y(N102) );
  INVX1 U135 ( .A(N222), .Y(n56) );
  OAI21X1 U136 ( .A(n2168), .B(n57), .C(reset_n), .Y(N101) );
  INVX1 U137 ( .A(N221), .Y(n57) );
  OAI21X1 U138 ( .A(n2168), .B(n58), .C(reset_n), .Y(N100) );
  INVX1 U139 ( .A(N220), .Y(n58) );
  NAND3X1 U140 ( .A(N129), .B(cs), .C(we), .Y(n24) );
  MUX2X1 U141 ( .B(core_block[1023]), .A(n2166), .S(n2222), .Y(n59) );
  INVX2 U142 ( .A(n59), .Y(n2106) );
  MUX2X1 U143 ( .B(core_block[1022]), .A(n2164), .S(n2222), .Y(n60) );
  INVX2 U144 ( .A(n60), .Y(n2105) );
  MUX2X1 U145 ( .B(core_block[1021]), .A(n2162), .S(n2222), .Y(n61) );
  INVX2 U146 ( .A(n61), .Y(n2104) );
  MUX2X1 U147 ( .B(core_block[1020]), .A(n2160), .S(n2222), .Y(n62) );
  INVX2 U148 ( .A(n62), .Y(n2103) );
  MUX2X1 U149 ( .B(core_block[1019]), .A(n2158), .S(n2222), .Y(n63) );
  INVX2 U150 ( .A(n63), .Y(n2102) );
  MUX2X1 U151 ( .B(core_block[1018]), .A(n2156), .S(n2222), .Y(n64) );
  INVX2 U152 ( .A(n64), .Y(n2101) );
  MUX2X1 U153 ( .B(core_block[1017]), .A(n2154), .S(n2222), .Y(n65) );
  INVX2 U154 ( .A(n65), .Y(n2100) );
  MUX2X1 U155 ( .B(core_block[1016]), .A(n2152), .S(n2222), .Y(n66) );
  INVX2 U156 ( .A(n66), .Y(n2099) );
  MUX2X1 U157 ( .B(core_block[1015]), .A(n2150), .S(n2222), .Y(n67) );
  INVX2 U158 ( .A(n67), .Y(n2098) );
  MUX2X1 U159 ( .B(core_block[1014]), .A(n2148), .S(n2222), .Y(n68) );
  INVX2 U160 ( .A(n68), .Y(n2097) );
  MUX2X1 U161 ( .B(core_block[1013]), .A(n2146), .S(n2222), .Y(n69) );
  INVX2 U162 ( .A(n69), .Y(n2096) );
  MUX2X1 U163 ( .B(core_block[1012]), .A(n2144), .S(n2222), .Y(n70) );
  INVX2 U164 ( .A(n70), .Y(n2095) );
  MUX2X1 U165 ( .B(core_block[1011]), .A(n2142), .S(n2222), .Y(n71) );
  INVX2 U166 ( .A(n71), .Y(n2094) );
  MUX2X1 U167 ( .B(core_block[1010]), .A(n2140), .S(n2222), .Y(n72) );
  INVX2 U168 ( .A(n72), .Y(n2093) );
  MUX2X1 U169 ( .B(core_block[1009]), .A(n2138), .S(n2222), .Y(n73) );
  INVX2 U170 ( .A(n73), .Y(n2092) );
  MUX2X1 U171 ( .B(core_block[1008]), .A(n2136), .S(n2222), .Y(n74) );
  INVX2 U172 ( .A(n74), .Y(n2091) );
  MUX2X1 U173 ( .B(core_block[1007]), .A(n2134), .S(n2222), .Y(n75) );
  INVX2 U174 ( .A(n75), .Y(n2090) );
  MUX2X1 U175 ( .B(core_block[1006]), .A(n2132), .S(n2222), .Y(n76) );
  INVX2 U176 ( .A(n76), .Y(n2089) );
  MUX2X1 U177 ( .B(core_block[1005]), .A(n2130), .S(n2222), .Y(n77) );
  INVX2 U178 ( .A(n77), .Y(n2088) );
  MUX2X1 U179 ( .B(core_block[1004]), .A(n2128), .S(n2222), .Y(n78) );
  INVX2 U180 ( .A(n78), .Y(n2087) );
  MUX2X1 U181 ( .B(core_block[1003]), .A(n2126), .S(n2222), .Y(n79) );
  INVX2 U182 ( .A(n79), .Y(n2086) );
  MUX2X1 U183 ( .B(core_block[1002]), .A(n2124), .S(n2222), .Y(n80) );
  INVX2 U184 ( .A(n80), .Y(n2085) );
  MUX2X1 U185 ( .B(core_block[1001]), .A(n2122), .S(n2222), .Y(n81) );
  INVX2 U186 ( .A(n81), .Y(n2084) );
  MUX2X1 U187 ( .B(core_block[1000]), .A(n2120), .S(n2222), .Y(n82) );
  INVX2 U188 ( .A(n82), .Y(n2083) );
  MUX2X1 U189 ( .B(core_block[999]), .A(n2118), .S(n2222), .Y(n83) );
  INVX2 U190 ( .A(n83), .Y(n2082) );
  MUX2X1 U191 ( .B(core_block[998]), .A(n2116), .S(n2222), .Y(n84) );
  INVX2 U192 ( .A(n84), .Y(n2081) );
  MUX2X1 U193 ( .B(core_block[997]), .A(n2114), .S(n2222), .Y(n85) );
  INVX2 U194 ( .A(n85), .Y(n2080) );
  MUX2X1 U195 ( .B(core_block[996]), .A(n2112), .S(n2222), .Y(n86) );
  INVX2 U196 ( .A(n86), .Y(n2079) );
  MUX2X1 U197 ( .B(core_block[995]), .A(n2110), .S(n2222), .Y(n87) );
  INVX2 U198 ( .A(n87), .Y(n2078) );
  MUX2X1 U199 ( .B(core_block[994]), .A(n2108), .S(n2222), .Y(n88) );
  INVX2 U200 ( .A(n88), .Y(n2077) );
  MUX2X1 U201 ( .B(core_block[993]), .A(n2172), .S(n2222), .Y(n89) );
  INVX2 U202 ( .A(n89), .Y(n2076) );
  MUX2X1 U203 ( .B(core_block[992]), .A(n2170), .S(n2222), .Y(n90) );
  INVX2 U204 ( .A(n90), .Y(n2075) );
  MUX2X1 U205 ( .B(core_block[991]), .A(n2166), .S(n2220), .Y(n91) );
  INVX2 U206 ( .A(n91), .Y(n2074) );
  MUX2X1 U207 ( .B(core_block[990]), .A(n2164), .S(n2220), .Y(n92) );
  INVX2 U208 ( .A(n92), .Y(n2073) );
  MUX2X1 U209 ( .B(core_block[989]), .A(n2162), .S(n2220), .Y(n93) );
  INVX2 U210 ( .A(n93), .Y(n2072) );
  MUX2X1 U211 ( .B(core_block[988]), .A(n2160), .S(n2220), .Y(n94) );
  INVX2 U212 ( .A(n94), .Y(n2071) );
  MUX2X1 U213 ( .B(core_block[987]), .A(n2158), .S(n2220), .Y(n95) );
  INVX2 U214 ( .A(n95), .Y(n2070) );
  MUX2X1 U215 ( .B(core_block[986]), .A(n2156), .S(n2220), .Y(n96) );
  INVX2 U216 ( .A(n96), .Y(n2069) );
  MUX2X1 U217 ( .B(core_block[985]), .A(n2154), .S(n2220), .Y(n97) );
  INVX2 U218 ( .A(n97), .Y(n2068) );
  MUX2X1 U219 ( .B(core_block[984]), .A(n2152), .S(n2220), .Y(n98) );
  INVX2 U220 ( .A(n98), .Y(n2067) );
  MUX2X1 U221 ( .B(core_block[983]), .A(n2150), .S(n2220), .Y(n99) );
  INVX2 U222 ( .A(n99), .Y(n2066) );
  MUX2X1 U223 ( .B(core_block[982]), .A(n2148), .S(n2220), .Y(n100) );
  INVX2 U224 ( .A(n100), .Y(n2065) );
  MUX2X1 U225 ( .B(core_block[981]), .A(n2146), .S(n2220), .Y(n101) );
  INVX2 U226 ( .A(n101), .Y(n2064) );
  MUX2X1 U227 ( .B(core_block[980]), .A(n2144), .S(n2220), .Y(n102) );
  INVX2 U228 ( .A(n102), .Y(n2063) );
  MUX2X1 U229 ( .B(core_block[979]), .A(n2142), .S(n2220), .Y(n103) );
  INVX2 U230 ( .A(n103), .Y(n2062) );
  MUX2X1 U231 ( .B(core_block[978]), .A(n2140), .S(n2220), .Y(n104) );
  INVX2 U232 ( .A(n104), .Y(n2061) );
  MUX2X1 U233 ( .B(core_block[977]), .A(n2138), .S(n2220), .Y(n105) );
  INVX2 U234 ( .A(n105), .Y(n2060) );
  MUX2X1 U235 ( .B(core_block[976]), .A(n2136), .S(n2220), .Y(n106) );
  INVX2 U236 ( .A(n106), .Y(n2059) );
  MUX2X1 U237 ( .B(core_block[975]), .A(n2134), .S(n2220), .Y(n107) );
  INVX2 U238 ( .A(n107), .Y(n2058) );
  MUX2X1 U239 ( .B(core_block[974]), .A(n2132), .S(n2220), .Y(n108) );
  INVX2 U240 ( .A(n108), .Y(n2057) );
  MUX2X1 U241 ( .B(core_block[973]), .A(n2130), .S(n2220), .Y(n109) );
  INVX2 U242 ( .A(n109), .Y(n2056) );
  MUX2X1 U243 ( .B(core_block[972]), .A(n2128), .S(n2220), .Y(n110) );
  INVX2 U244 ( .A(n110), .Y(n2055) );
  MUX2X1 U245 ( .B(core_block[971]), .A(n2126), .S(n2220), .Y(n111) );
  INVX2 U246 ( .A(n111), .Y(n2054) );
  MUX2X1 U247 ( .B(core_block[970]), .A(n2124), .S(n2220), .Y(n112) );
  INVX2 U248 ( .A(n112), .Y(n2053) );
  MUX2X1 U249 ( .B(core_block[969]), .A(n2122), .S(n2220), .Y(n113) );
  INVX2 U250 ( .A(n113), .Y(n2052) );
  MUX2X1 U251 ( .B(core_block[968]), .A(n2120), .S(n2220), .Y(n114) );
  INVX2 U252 ( .A(n114), .Y(n2051) );
  MUX2X1 U253 ( .B(core_block[967]), .A(n2118), .S(n2220), .Y(n115) );
  INVX2 U254 ( .A(n115), .Y(n2050) );
  MUX2X1 U255 ( .B(core_block[966]), .A(n2116), .S(n2220), .Y(n116) );
  INVX2 U256 ( .A(n116), .Y(n2049) );
  MUX2X1 U257 ( .B(core_block[965]), .A(n2114), .S(n2220), .Y(n117) );
  INVX2 U258 ( .A(n117), .Y(n2048) );
  MUX2X1 U259 ( .B(core_block[964]), .A(n2112), .S(n2220), .Y(n118) );
  INVX2 U260 ( .A(n118), .Y(n2047) );
  MUX2X1 U261 ( .B(core_block[963]), .A(n2110), .S(n2220), .Y(n119) );
  INVX2 U262 ( .A(n119), .Y(n2046) );
  MUX2X1 U263 ( .B(core_block[962]), .A(n2108), .S(n2220), .Y(n120) );
  INVX2 U264 ( .A(n120), .Y(n2045) );
  MUX2X1 U265 ( .B(core_block[961]), .A(n2172), .S(n2220), .Y(n121) );
  INVX2 U266 ( .A(n121), .Y(n2044) );
  MUX2X1 U267 ( .B(core_block[960]), .A(n2170), .S(n2220), .Y(n122) );
  INVX2 U268 ( .A(n122), .Y(n2043) );
  MUX2X1 U269 ( .B(core_block[959]), .A(n2166), .S(n2218), .Y(n123) );
  INVX2 U270 ( .A(n123), .Y(n2042) );
  MUX2X1 U271 ( .B(core_block[958]), .A(n2164), .S(n2218), .Y(n124) );
  INVX2 U272 ( .A(n124), .Y(n2041) );
  MUX2X1 U273 ( .B(core_block[957]), .A(n2162), .S(n2218), .Y(n125) );
  INVX2 U274 ( .A(n125), .Y(n2040) );
  MUX2X1 U275 ( .B(core_block[956]), .A(n2160), .S(n2218), .Y(n126) );
  INVX2 U276 ( .A(n126), .Y(n2039) );
  MUX2X1 U277 ( .B(core_block[955]), .A(n2158), .S(n2218), .Y(n127) );
  INVX2 U278 ( .A(n127), .Y(n2038) );
  MUX2X1 U279 ( .B(core_block[954]), .A(n2156), .S(n2218), .Y(n128) );
  INVX2 U280 ( .A(n128), .Y(n2037) );
  MUX2X1 U281 ( .B(core_block[953]), .A(n2154), .S(n2218), .Y(n129) );
  INVX2 U282 ( .A(n129), .Y(n2036) );
  MUX2X1 U283 ( .B(core_block[952]), .A(n2152), .S(n2218), .Y(n130) );
  INVX2 U284 ( .A(n130), .Y(n2035) );
  MUX2X1 U285 ( .B(core_block[951]), .A(n2150), .S(n2218), .Y(n131) );
  INVX2 U286 ( .A(n131), .Y(n2034) );
  MUX2X1 U287 ( .B(core_block[950]), .A(n2148), .S(n2218), .Y(n132) );
  INVX2 U288 ( .A(n132), .Y(n2033) );
  MUX2X1 U289 ( .B(core_block[949]), .A(n2146), .S(n2218), .Y(n133) );
  INVX2 U290 ( .A(n133), .Y(n2032) );
  MUX2X1 U291 ( .B(core_block[948]), .A(n2144), .S(n2218), .Y(n134) );
  INVX2 U292 ( .A(n134), .Y(n2031) );
  MUX2X1 U293 ( .B(core_block[947]), .A(n2142), .S(n2218), .Y(n135) );
  INVX2 U294 ( .A(n135), .Y(n2030) );
  MUX2X1 U295 ( .B(core_block[946]), .A(n2140), .S(n2218), .Y(n136) );
  INVX2 U296 ( .A(n136), .Y(n2029) );
  MUX2X1 U297 ( .B(core_block[945]), .A(n2138), .S(n2218), .Y(n137) );
  INVX2 U298 ( .A(n137), .Y(n2028) );
  MUX2X1 U299 ( .B(core_block[944]), .A(n2136), .S(n2218), .Y(n138) );
  INVX2 U300 ( .A(n138), .Y(n2027) );
  MUX2X1 U301 ( .B(core_block[943]), .A(n2134), .S(n2218), .Y(n139) );
  INVX2 U302 ( .A(n139), .Y(n2026) );
  MUX2X1 U303 ( .B(core_block[942]), .A(n2132), .S(n2218), .Y(n140) );
  INVX2 U304 ( .A(n140), .Y(n2025) );
  MUX2X1 U305 ( .B(core_block[941]), .A(n2130), .S(n2218), .Y(n141) );
  INVX2 U306 ( .A(n141), .Y(n2024) );
  MUX2X1 U307 ( .B(core_block[940]), .A(n2128), .S(n2218), .Y(n142) );
  INVX2 U308 ( .A(n142), .Y(n2023) );
  MUX2X1 U309 ( .B(core_block[939]), .A(n2126), .S(n2218), .Y(n143) );
  INVX2 U310 ( .A(n143), .Y(n2022) );
  MUX2X1 U311 ( .B(core_block[938]), .A(n2124), .S(n2218), .Y(n144) );
  INVX2 U312 ( .A(n144), .Y(n2021) );
  MUX2X1 U313 ( .B(core_block[937]), .A(n2122), .S(n2218), .Y(n145) );
  INVX2 U314 ( .A(n145), .Y(n2020) );
  MUX2X1 U315 ( .B(core_block[936]), .A(n2120), .S(n2218), .Y(n146) );
  INVX2 U316 ( .A(n146), .Y(n2019) );
  MUX2X1 U317 ( .B(core_block[935]), .A(n2118), .S(n2218), .Y(n147) );
  INVX2 U318 ( .A(n147), .Y(n2018) );
  MUX2X1 U319 ( .B(core_block[934]), .A(n2116), .S(n2218), .Y(n148) );
  INVX2 U320 ( .A(n148), .Y(n2017) );
  MUX2X1 U321 ( .B(core_block[933]), .A(n2114), .S(n2218), .Y(n149) );
  INVX2 U322 ( .A(n149), .Y(n2016) );
  MUX2X1 U323 ( .B(core_block[932]), .A(n2112), .S(n2218), .Y(n150) );
  INVX2 U324 ( .A(n150), .Y(n2015) );
  MUX2X1 U325 ( .B(core_block[931]), .A(n2110), .S(n2218), .Y(n151) );
  INVX2 U326 ( .A(n151), .Y(n2014) );
  MUX2X1 U327 ( .B(core_block[930]), .A(n2108), .S(n2218), .Y(n152) );
  INVX2 U328 ( .A(n152), .Y(n2013) );
  MUX2X1 U329 ( .B(core_block[929]), .A(n2172), .S(n2218), .Y(n153) );
  INVX2 U330 ( .A(n153), .Y(n2012) );
  MUX2X1 U331 ( .B(core_block[928]), .A(n2170), .S(n2218), .Y(n154) );
  INVX2 U332 ( .A(n154), .Y(n2011) );
  MUX2X1 U333 ( .B(core_block[927]), .A(n2166), .S(n2216), .Y(n155) );
  INVX2 U334 ( .A(n155), .Y(n2010) );
  MUX2X1 U335 ( .B(core_block[926]), .A(n2164), .S(n2216), .Y(n156) );
  INVX2 U336 ( .A(n156), .Y(n2009) );
  MUX2X1 U337 ( .B(core_block[925]), .A(n2162), .S(n2216), .Y(n157) );
  INVX2 U338 ( .A(n157), .Y(n2008) );
  MUX2X1 U339 ( .B(core_block[924]), .A(n2160), .S(n2216), .Y(n158) );
  INVX2 U340 ( .A(n158), .Y(n2007) );
  MUX2X1 U341 ( .B(core_block[923]), .A(n2158), .S(n2216), .Y(n159) );
  INVX2 U342 ( .A(n159), .Y(n2006) );
  MUX2X1 U343 ( .B(core_block[922]), .A(n2156), .S(n2216), .Y(n160) );
  INVX2 U344 ( .A(n160), .Y(n2005) );
  MUX2X1 U345 ( .B(core_block[921]), .A(n2154), .S(n2216), .Y(n161) );
  INVX2 U346 ( .A(n161), .Y(n2004) );
  MUX2X1 U347 ( .B(core_block[920]), .A(n2152), .S(n2216), .Y(n162) );
  INVX2 U348 ( .A(n162), .Y(n2003) );
  MUX2X1 U349 ( .B(core_block[919]), .A(n2150), .S(n2216), .Y(n163) );
  INVX2 U350 ( .A(n163), .Y(n2002) );
  MUX2X1 U351 ( .B(core_block[918]), .A(n2148), .S(n2216), .Y(n164) );
  INVX2 U352 ( .A(n164), .Y(n2001) );
  MUX2X1 U353 ( .B(core_block[917]), .A(n2146), .S(n2216), .Y(n165) );
  INVX2 U354 ( .A(n165), .Y(n2000) );
  MUX2X1 U355 ( .B(core_block[916]), .A(n2144), .S(n2216), .Y(n166) );
  INVX2 U356 ( .A(n166), .Y(n1999) );
  MUX2X1 U357 ( .B(core_block[915]), .A(n2142), .S(n2216), .Y(n167) );
  INVX2 U358 ( .A(n167), .Y(n1998) );
  MUX2X1 U359 ( .B(core_block[914]), .A(n2140), .S(n2216), .Y(n168) );
  INVX2 U360 ( .A(n168), .Y(n1997) );
  MUX2X1 U361 ( .B(core_block[913]), .A(n2138), .S(n2216), .Y(n169) );
  INVX2 U362 ( .A(n169), .Y(n1996) );
  MUX2X1 U363 ( .B(core_block[912]), .A(n2136), .S(n2216), .Y(n170) );
  INVX2 U364 ( .A(n170), .Y(n1995) );
  MUX2X1 U365 ( .B(core_block[911]), .A(n2134), .S(n2216), .Y(n171) );
  INVX2 U366 ( .A(n171), .Y(n1994) );
  MUX2X1 U367 ( .B(core_block[910]), .A(n2132), .S(n2216), .Y(n172) );
  INVX2 U368 ( .A(n172), .Y(n1993) );
  MUX2X1 U369 ( .B(core_block[909]), .A(n2130), .S(n2216), .Y(n173) );
  INVX2 U370 ( .A(n173), .Y(n1992) );
  MUX2X1 U371 ( .B(core_block[908]), .A(n2128), .S(n2216), .Y(n174) );
  INVX2 U372 ( .A(n174), .Y(n1991) );
  MUX2X1 U373 ( .B(core_block[907]), .A(n2126), .S(n2216), .Y(n175) );
  INVX2 U374 ( .A(n175), .Y(n1990) );
  MUX2X1 U375 ( .B(core_block[906]), .A(n2124), .S(n2216), .Y(n176) );
  INVX2 U376 ( .A(n176), .Y(n1989) );
  MUX2X1 U377 ( .B(core_block[905]), .A(n2122), .S(n2216), .Y(n177) );
  INVX2 U378 ( .A(n177), .Y(n1988) );
  MUX2X1 U379 ( .B(core_block[904]), .A(n2120), .S(n2216), .Y(n178) );
  INVX2 U380 ( .A(n178), .Y(n1987) );
  MUX2X1 U381 ( .B(core_block[903]), .A(n2118), .S(n2216), .Y(n179) );
  INVX2 U382 ( .A(n179), .Y(n1986) );
  MUX2X1 U383 ( .B(core_block[902]), .A(n2116), .S(n2216), .Y(n180) );
  INVX2 U384 ( .A(n180), .Y(n1985) );
  MUX2X1 U385 ( .B(core_block[901]), .A(n2114), .S(n2216), .Y(n181) );
  INVX2 U386 ( .A(n181), .Y(n1984) );
  MUX2X1 U387 ( .B(core_block[900]), .A(n2112), .S(n2216), .Y(n182) );
  INVX2 U388 ( .A(n182), .Y(n1983) );
  MUX2X1 U389 ( .B(core_block[899]), .A(n2110), .S(n2216), .Y(n183) );
  INVX2 U390 ( .A(n183), .Y(n1982) );
  MUX2X1 U391 ( .B(core_block[898]), .A(n2108), .S(n2216), .Y(n184) );
  INVX2 U392 ( .A(n184), .Y(n1981) );
  MUX2X1 U393 ( .B(core_block[897]), .A(n2172), .S(n2216), .Y(n185) );
  INVX2 U394 ( .A(n185), .Y(n1980) );
  MUX2X1 U395 ( .B(core_block[896]), .A(n2170), .S(n2216), .Y(n186) );
  INVX2 U396 ( .A(n186), .Y(n1979) );
  MUX2X1 U397 ( .B(core_block[895]), .A(n2166), .S(n2214), .Y(n187) );
  INVX2 U398 ( .A(n187), .Y(n1978) );
  MUX2X1 U399 ( .B(core_block[894]), .A(n2164), .S(n2214), .Y(n188) );
  INVX2 U400 ( .A(n188), .Y(n1977) );
  MUX2X1 U401 ( .B(core_block[893]), .A(n2162), .S(n2214), .Y(n189) );
  INVX2 U402 ( .A(n189), .Y(n1976) );
  MUX2X1 U403 ( .B(core_block[892]), .A(n2160), .S(n2214), .Y(n190) );
  INVX2 U404 ( .A(n190), .Y(n1975) );
  MUX2X1 U405 ( .B(core_block[891]), .A(n2158), .S(n2214), .Y(n191) );
  INVX2 U406 ( .A(n191), .Y(n1974) );
  MUX2X1 U407 ( .B(core_block[890]), .A(n2156), .S(n2214), .Y(n192) );
  INVX2 U408 ( .A(n192), .Y(n1973) );
  MUX2X1 U409 ( .B(core_block[889]), .A(n2154), .S(n2214), .Y(n193) );
  INVX2 U410 ( .A(n193), .Y(n1972) );
  MUX2X1 U411 ( .B(core_block[888]), .A(n2152), .S(n2214), .Y(n194) );
  INVX2 U412 ( .A(n194), .Y(n1971) );
  MUX2X1 U413 ( .B(core_block[887]), .A(n2150), .S(n2214), .Y(n195) );
  INVX2 U414 ( .A(n195), .Y(n1970) );
  MUX2X1 U415 ( .B(core_block[886]), .A(n2148), .S(n2214), .Y(n196) );
  INVX2 U416 ( .A(n196), .Y(n1969) );
  MUX2X1 U417 ( .B(core_block[885]), .A(n2146), .S(n2214), .Y(n197) );
  INVX2 U418 ( .A(n197), .Y(n1968) );
  MUX2X1 U419 ( .B(core_block[884]), .A(n2144), .S(n2214), .Y(n198) );
  INVX2 U420 ( .A(n198), .Y(n1967) );
  MUX2X1 U421 ( .B(core_block[883]), .A(n2142), .S(n2214), .Y(n199) );
  INVX2 U422 ( .A(n199), .Y(n1966) );
  MUX2X1 U423 ( .B(core_block[882]), .A(n2140), .S(n2214), .Y(n200) );
  INVX2 U424 ( .A(n200), .Y(n1965) );
  MUX2X1 U425 ( .B(core_block[881]), .A(n2138), .S(n2214), .Y(n201) );
  INVX2 U426 ( .A(n201), .Y(n1964) );
  MUX2X1 U427 ( .B(core_block[880]), .A(n2136), .S(n2214), .Y(n202) );
  INVX2 U428 ( .A(n202), .Y(n1963) );
  MUX2X1 U429 ( .B(core_block[879]), .A(n2134), .S(n2214), .Y(n203) );
  INVX2 U430 ( .A(n203), .Y(n1962) );
  MUX2X1 U431 ( .B(core_block[878]), .A(n2132), .S(n2214), .Y(n204) );
  INVX2 U432 ( .A(n204), .Y(n1961) );
  MUX2X1 U433 ( .B(core_block[877]), .A(n2130), .S(n2214), .Y(n205) );
  INVX2 U434 ( .A(n205), .Y(n1960) );
  MUX2X1 U435 ( .B(core_block[876]), .A(n2128), .S(n2214), .Y(n206) );
  INVX2 U436 ( .A(n206), .Y(n1959) );
  MUX2X1 U437 ( .B(core_block[875]), .A(n2126), .S(n2214), .Y(n207) );
  INVX2 U438 ( .A(n207), .Y(n1958) );
  MUX2X1 U439 ( .B(core_block[874]), .A(n2124), .S(n2214), .Y(n208) );
  INVX2 U440 ( .A(n208), .Y(n1957) );
  MUX2X1 U441 ( .B(core_block[873]), .A(n2122), .S(n2214), .Y(n209) );
  INVX2 U442 ( .A(n209), .Y(n1956) );
  MUX2X1 U443 ( .B(core_block[872]), .A(n2120), .S(n2214), .Y(n210) );
  INVX2 U444 ( .A(n210), .Y(n1955) );
  MUX2X1 U445 ( .B(core_block[871]), .A(n2118), .S(n2214), .Y(n211) );
  INVX2 U446 ( .A(n211), .Y(n1954) );
  MUX2X1 U447 ( .B(core_block[870]), .A(n2116), .S(n2214), .Y(n212) );
  INVX2 U448 ( .A(n212), .Y(n1953) );
  MUX2X1 U449 ( .B(core_block[869]), .A(n2114), .S(n2214), .Y(n213) );
  INVX2 U450 ( .A(n213), .Y(n1952) );
  MUX2X1 U451 ( .B(core_block[868]), .A(n2112), .S(n2214), .Y(n214) );
  INVX2 U452 ( .A(n214), .Y(n1951) );
  MUX2X1 U453 ( .B(core_block[867]), .A(n2110), .S(n2214), .Y(n215) );
  INVX2 U454 ( .A(n215), .Y(n1950) );
  MUX2X1 U455 ( .B(core_block[866]), .A(n2108), .S(n2214), .Y(n216) );
  INVX2 U456 ( .A(n216), .Y(n1949) );
  MUX2X1 U457 ( .B(core_block[865]), .A(n2172), .S(n2214), .Y(n217) );
  INVX2 U458 ( .A(n217), .Y(n1948) );
  MUX2X1 U459 ( .B(core_block[864]), .A(n2170), .S(n2214), .Y(n218) );
  INVX2 U460 ( .A(n218), .Y(n1947) );
  MUX2X1 U461 ( .B(core_block[863]), .A(n2166), .S(n2212), .Y(n219) );
  INVX2 U462 ( .A(n219), .Y(n1946) );
  MUX2X1 U463 ( .B(core_block[862]), .A(n2164), .S(n2212), .Y(n220) );
  INVX2 U464 ( .A(n220), .Y(n1945) );
  MUX2X1 U465 ( .B(core_block[861]), .A(n2162), .S(n2212), .Y(n221) );
  INVX2 U466 ( .A(n221), .Y(n1944) );
  MUX2X1 U467 ( .B(core_block[860]), .A(n2160), .S(n2212), .Y(n222) );
  INVX2 U468 ( .A(n222), .Y(n1943) );
  MUX2X1 U469 ( .B(core_block[859]), .A(n2158), .S(n2212), .Y(n223) );
  INVX2 U470 ( .A(n223), .Y(n1942) );
  MUX2X1 U471 ( .B(core_block[858]), .A(n2156), .S(n2212), .Y(n224) );
  INVX2 U472 ( .A(n224), .Y(n1941) );
  MUX2X1 U473 ( .B(core_block[857]), .A(n2154), .S(n2212), .Y(n225) );
  INVX2 U474 ( .A(n225), .Y(n1940) );
  MUX2X1 U475 ( .B(core_block[856]), .A(n2152), .S(n2212), .Y(n226) );
  INVX2 U476 ( .A(n226), .Y(n1939) );
  MUX2X1 U477 ( .B(core_block[855]), .A(n2150), .S(n2212), .Y(n227) );
  INVX2 U478 ( .A(n227), .Y(n1938) );
  MUX2X1 U479 ( .B(core_block[854]), .A(n2148), .S(n2212), .Y(n228) );
  INVX2 U480 ( .A(n228), .Y(n1937) );
  MUX2X1 U481 ( .B(core_block[853]), .A(n2146), .S(n2212), .Y(n229) );
  INVX2 U482 ( .A(n229), .Y(n1936) );
  MUX2X1 U483 ( .B(core_block[852]), .A(n2144), .S(n2212), .Y(n230) );
  INVX2 U484 ( .A(n230), .Y(n1935) );
  MUX2X1 U485 ( .B(core_block[851]), .A(n2142), .S(n2212), .Y(n231) );
  INVX2 U486 ( .A(n231), .Y(n1934) );
  MUX2X1 U487 ( .B(core_block[850]), .A(n2140), .S(n2212), .Y(n232) );
  INVX2 U488 ( .A(n232), .Y(n1933) );
  MUX2X1 U489 ( .B(core_block[849]), .A(n2138), .S(n2212), .Y(n233) );
  INVX2 U490 ( .A(n233), .Y(n1932) );
  MUX2X1 U491 ( .B(core_block[848]), .A(n2136), .S(n2212), .Y(n234) );
  INVX2 U492 ( .A(n234), .Y(n1931) );
  MUX2X1 U493 ( .B(core_block[847]), .A(n2134), .S(n2212), .Y(n235) );
  INVX2 U494 ( .A(n235), .Y(n1930) );
  MUX2X1 U495 ( .B(core_block[846]), .A(n2132), .S(n2212), .Y(n236) );
  INVX2 U496 ( .A(n236), .Y(n1929) );
  MUX2X1 U497 ( .B(core_block[845]), .A(n2130), .S(n2212), .Y(n237) );
  INVX2 U498 ( .A(n237), .Y(n1928) );
  MUX2X1 U499 ( .B(core_block[844]), .A(n2128), .S(n2212), .Y(n238) );
  INVX2 U500 ( .A(n238), .Y(n1927) );
  MUX2X1 U501 ( .B(core_block[843]), .A(n2126), .S(n2212), .Y(n239) );
  INVX2 U502 ( .A(n239), .Y(n1926) );
  MUX2X1 U503 ( .B(core_block[842]), .A(n2124), .S(n2212), .Y(n240) );
  INVX2 U504 ( .A(n240), .Y(n1925) );
  MUX2X1 U505 ( .B(core_block[841]), .A(n2122), .S(n2212), .Y(n241) );
  INVX2 U506 ( .A(n241), .Y(n1924) );
  MUX2X1 U507 ( .B(core_block[840]), .A(n2120), .S(n2212), .Y(n242) );
  INVX2 U508 ( .A(n242), .Y(n1923) );
  MUX2X1 U509 ( .B(core_block[839]), .A(n2118), .S(n2212), .Y(n243) );
  INVX2 U510 ( .A(n243), .Y(n1922) );
  MUX2X1 U511 ( .B(core_block[838]), .A(n2116), .S(n2212), .Y(n244) );
  INVX2 U512 ( .A(n244), .Y(n1921) );
  MUX2X1 U513 ( .B(core_block[837]), .A(n2114), .S(n2212), .Y(n245) );
  INVX2 U514 ( .A(n245), .Y(n1920) );
  MUX2X1 U515 ( .B(core_block[836]), .A(n2112), .S(n2212), .Y(n246) );
  INVX2 U516 ( .A(n246), .Y(n1919) );
  MUX2X1 U517 ( .B(core_block[835]), .A(n2110), .S(n2212), .Y(n247) );
  INVX2 U518 ( .A(n247), .Y(n1918) );
  MUX2X1 U519 ( .B(core_block[834]), .A(n2108), .S(n2212), .Y(n248) );
  INVX2 U520 ( .A(n248), .Y(n1917) );
  MUX2X1 U521 ( .B(core_block[833]), .A(n2172), .S(n2212), .Y(n249) );
  INVX2 U522 ( .A(n249), .Y(n1916) );
  MUX2X1 U523 ( .B(core_block[832]), .A(n2170), .S(n2212), .Y(n250) );
  INVX2 U524 ( .A(n250), .Y(n1915) );
  MUX2X1 U525 ( .B(core_block[831]), .A(n2166), .S(n2210), .Y(n251) );
  INVX2 U526 ( .A(n251), .Y(n1914) );
  MUX2X1 U527 ( .B(core_block[830]), .A(n2164), .S(n2210), .Y(n252) );
  INVX2 U528 ( .A(n252), .Y(n1913) );
  MUX2X1 U529 ( .B(core_block[829]), .A(n2162), .S(n2210), .Y(n253) );
  INVX2 U530 ( .A(n253), .Y(n1912) );
  MUX2X1 U531 ( .B(core_block[828]), .A(n2160), .S(n2210), .Y(n254) );
  INVX2 U532 ( .A(n254), .Y(n1911) );
  MUX2X1 U533 ( .B(core_block[827]), .A(n2158), .S(n2210), .Y(n255) );
  INVX2 U534 ( .A(n255), .Y(n1910) );
  MUX2X1 U535 ( .B(core_block[826]), .A(n2156), .S(n2210), .Y(n256) );
  INVX2 U536 ( .A(n256), .Y(n1909) );
  MUX2X1 U537 ( .B(core_block[825]), .A(n2154), .S(n2210), .Y(n257) );
  INVX2 U538 ( .A(n257), .Y(n1908) );
  MUX2X1 U539 ( .B(core_block[824]), .A(n2152), .S(n2210), .Y(n258) );
  INVX2 U540 ( .A(n258), .Y(n1907) );
  MUX2X1 U541 ( .B(core_block[823]), .A(n2150), .S(n2210), .Y(n259) );
  INVX2 U542 ( .A(n259), .Y(n1906) );
  MUX2X1 U543 ( .B(core_block[822]), .A(n2148), .S(n2210), .Y(n260) );
  INVX2 U544 ( .A(n260), .Y(n1905) );
  MUX2X1 U545 ( .B(core_block[821]), .A(n2146), .S(n2210), .Y(n261) );
  INVX2 U546 ( .A(n261), .Y(n1904) );
  MUX2X1 U547 ( .B(core_block[820]), .A(n2144), .S(n2210), .Y(n262) );
  INVX2 U548 ( .A(n262), .Y(n1903) );
  MUX2X1 U549 ( .B(core_block[819]), .A(n2142), .S(n2210), .Y(n263) );
  INVX2 U550 ( .A(n263), .Y(n1902) );
  MUX2X1 U551 ( .B(core_block[818]), .A(n2140), .S(n2210), .Y(n264) );
  INVX2 U552 ( .A(n264), .Y(n1901) );
  MUX2X1 U553 ( .B(core_block[817]), .A(n2138), .S(n2210), .Y(n265) );
  INVX2 U554 ( .A(n265), .Y(n1900) );
  MUX2X1 U555 ( .B(core_block[816]), .A(n2136), .S(n2210), .Y(n266) );
  INVX2 U556 ( .A(n266), .Y(n1899) );
  MUX2X1 U557 ( .B(core_block[815]), .A(n2134), .S(n2210), .Y(n267) );
  INVX2 U558 ( .A(n267), .Y(n1898) );
  MUX2X1 U559 ( .B(core_block[814]), .A(n2132), .S(n2210), .Y(n268) );
  INVX2 U560 ( .A(n268), .Y(n1897) );
  MUX2X1 U561 ( .B(core_block[813]), .A(n2130), .S(n2210), .Y(n269) );
  INVX2 U562 ( .A(n269), .Y(n1896) );
  MUX2X1 U563 ( .B(core_block[812]), .A(n2128), .S(n2210), .Y(n270) );
  INVX2 U564 ( .A(n270), .Y(n1895) );
  MUX2X1 U565 ( .B(core_block[811]), .A(n2126), .S(n2210), .Y(n271) );
  INVX2 U566 ( .A(n271), .Y(n1894) );
  MUX2X1 U567 ( .B(core_block[810]), .A(n2124), .S(n2210), .Y(n272) );
  INVX2 U568 ( .A(n272), .Y(n1893) );
  MUX2X1 U569 ( .B(core_block[809]), .A(n2122), .S(n2210), .Y(n273) );
  INVX2 U570 ( .A(n273), .Y(n1892) );
  MUX2X1 U571 ( .B(core_block[808]), .A(n2120), .S(n2210), .Y(n274) );
  INVX2 U572 ( .A(n274), .Y(n1891) );
  MUX2X1 U573 ( .B(core_block[807]), .A(n2118), .S(n2210), .Y(n275) );
  INVX2 U574 ( .A(n275), .Y(n1890) );
  MUX2X1 U575 ( .B(core_block[806]), .A(n2116), .S(n2210), .Y(n276) );
  INVX2 U576 ( .A(n276), .Y(n1889) );
  MUX2X1 U577 ( .B(core_block[805]), .A(n2114), .S(n2210), .Y(n277) );
  INVX2 U578 ( .A(n277), .Y(n1888) );
  MUX2X1 U579 ( .B(core_block[804]), .A(n2112), .S(n2210), .Y(n278) );
  INVX2 U580 ( .A(n278), .Y(n1887) );
  MUX2X1 U581 ( .B(core_block[803]), .A(n2110), .S(n2210), .Y(n279) );
  INVX2 U582 ( .A(n279), .Y(n1886) );
  MUX2X1 U583 ( .B(core_block[802]), .A(n2108), .S(n2210), .Y(n280) );
  INVX2 U584 ( .A(n280), .Y(n1885) );
  MUX2X1 U585 ( .B(core_block[801]), .A(n2172), .S(n2210), .Y(n281) );
  INVX2 U586 ( .A(n281), .Y(n1884) );
  MUX2X1 U587 ( .B(core_block[800]), .A(n2170), .S(n2210), .Y(n282) );
  INVX2 U588 ( .A(n282), .Y(n1883) );
  MUX2X1 U589 ( .B(core_block[799]), .A(n2166), .S(n2208), .Y(n283) );
  INVX2 U590 ( .A(n283), .Y(n1882) );
  MUX2X1 U591 ( .B(core_block[798]), .A(n2164), .S(n2208), .Y(n284) );
  INVX2 U592 ( .A(n284), .Y(n1881) );
  MUX2X1 U593 ( .B(core_block[797]), .A(n2162), .S(n2208), .Y(n285) );
  INVX2 U594 ( .A(n285), .Y(n1880) );
  MUX2X1 U595 ( .B(core_block[796]), .A(n2160), .S(n2208), .Y(n286) );
  INVX2 U596 ( .A(n286), .Y(n1879) );
  MUX2X1 U597 ( .B(core_block[795]), .A(n2158), .S(n2208), .Y(n287) );
  INVX2 U598 ( .A(n287), .Y(n1878) );
  MUX2X1 U599 ( .B(core_block[794]), .A(n2156), .S(n2208), .Y(n288) );
  INVX2 U600 ( .A(n288), .Y(n1877) );
  MUX2X1 U601 ( .B(core_block[793]), .A(n2154), .S(n2208), .Y(n289) );
  INVX2 U602 ( .A(n289), .Y(n1876) );
  MUX2X1 U603 ( .B(core_block[792]), .A(n2152), .S(n2208), .Y(n290) );
  INVX2 U604 ( .A(n290), .Y(n1875) );
  MUX2X1 U605 ( .B(core_block[791]), .A(n2150), .S(n2208), .Y(n291) );
  INVX2 U606 ( .A(n291), .Y(n1874) );
  MUX2X1 U607 ( .B(core_block[790]), .A(n2148), .S(n2208), .Y(n292) );
  INVX2 U608 ( .A(n292), .Y(n1873) );
  MUX2X1 U609 ( .B(core_block[789]), .A(n2146), .S(n2208), .Y(n293) );
  INVX2 U610 ( .A(n293), .Y(n1872) );
  MUX2X1 U611 ( .B(core_block[788]), .A(n2144), .S(n2208), .Y(n294) );
  INVX2 U612 ( .A(n294), .Y(n1871) );
  MUX2X1 U613 ( .B(core_block[787]), .A(n2142), .S(n2208), .Y(n295) );
  INVX2 U614 ( .A(n295), .Y(n1870) );
  MUX2X1 U615 ( .B(core_block[786]), .A(n2140), .S(n2208), .Y(n296) );
  INVX2 U616 ( .A(n296), .Y(n1869) );
  MUX2X1 U617 ( .B(core_block[785]), .A(n2138), .S(n2208), .Y(n297) );
  INVX2 U618 ( .A(n297), .Y(n1868) );
  MUX2X1 U619 ( .B(core_block[784]), .A(n2136), .S(n2208), .Y(n298) );
  INVX2 U620 ( .A(n298), .Y(n1867) );
  MUX2X1 U621 ( .B(core_block[783]), .A(n2134), .S(n2208), .Y(n299) );
  INVX2 U622 ( .A(n299), .Y(n1866) );
  MUX2X1 U623 ( .B(core_block[782]), .A(n2132), .S(n2208), .Y(n300) );
  INVX2 U624 ( .A(n300), .Y(n1865) );
  MUX2X1 U625 ( .B(core_block[781]), .A(n2130), .S(n2208), .Y(n301) );
  INVX2 U626 ( .A(n301), .Y(n1864) );
  MUX2X1 U627 ( .B(core_block[780]), .A(n2128), .S(n2208), .Y(n302) );
  INVX2 U628 ( .A(n302), .Y(n1863) );
  MUX2X1 U629 ( .B(core_block[779]), .A(n2126), .S(n2208), .Y(n303) );
  INVX2 U630 ( .A(n303), .Y(n1862) );
  MUX2X1 U631 ( .B(core_block[778]), .A(n2124), .S(n2208), .Y(n304) );
  INVX2 U632 ( .A(n304), .Y(n1861) );
  MUX2X1 U633 ( .B(core_block[777]), .A(n2122), .S(n2208), .Y(n305) );
  INVX2 U634 ( .A(n305), .Y(n1860) );
  MUX2X1 U635 ( .B(core_block[776]), .A(n2120), .S(n2208), .Y(n306) );
  INVX2 U636 ( .A(n306), .Y(n1859) );
  MUX2X1 U637 ( .B(core_block[775]), .A(n2118), .S(n2208), .Y(n307) );
  INVX2 U638 ( .A(n307), .Y(n1858) );
  MUX2X1 U639 ( .B(core_block[774]), .A(n2116), .S(n2208), .Y(n308) );
  INVX2 U640 ( .A(n308), .Y(n1857) );
  MUX2X1 U641 ( .B(core_block[773]), .A(n2114), .S(n2208), .Y(n309) );
  INVX2 U642 ( .A(n309), .Y(n1856) );
  MUX2X1 U643 ( .B(core_block[772]), .A(n2112), .S(n2208), .Y(n310) );
  INVX2 U644 ( .A(n310), .Y(n1855) );
  MUX2X1 U645 ( .B(core_block[771]), .A(n2110), .S(n2208), .Y(n311) );
  INVX2 U646 ( .A(n311), .Y(n1854) );
  MUX2X1 U647 ( .B(core_block[770]), .A(n2108), .S(n2208), .Y(n312) );
  INVX2 U648 ( .A(n312), .Y(n1853) );
  MUX2X1 U649 ( .B(core_block[769]), .A(n2172), .S(n2208), .Y(n313) );
  INVX2 U650 ( .A(n313), .Y(n1852) );
  MUX2X1 U651 ( .B(core_block[768]), .A(n2170), .S(n2208), .Y(n314) );
  INVX2 U652 ( .A(n314), .Y(n1851) );
  MUX2X1 U653 ( .B(core_block[767]), .A(n2166), .S(n2206), .Y(n315) );
  INVX2 U654 ( .A(n315), .Y(n1850) );
  MUX2X1 U655 ( .B(core_block[766]), .A(n2164), .S(n2206), .Y(n316) );
  INVX2 U656 ( .A(n316), .Y(n1849) );
  MUX2X1 U657 ( .B(core_block[765]), .A(n2162), .S(n2206), .Y(n317) );
  INVX2 U658 ( .A(n317), .Y(n1848) );
  MUX2X1 U659 ( .B(core_block[764]), .A(n2160), .S(n2206), .Y(n318) );
  INVX2 U660 ( .A(n318), .Y(n1847) );
  MUX2X1 U661 ( .B(core_block[763]), .A(n2158), .S(n2206), .Y(n319) );
  INVX2 U662 ( .A(n319), .Y(n1846) );
  MUX2X1 U663 ( .B(core_block[762]), .A(n2156), .S(n2206), .Y(n320) );
  INVX2 U664 ( .A(n320), .Y(n1845) );
  MUX2X1 U665 ( .B(core_block[761]), .A(n2154), .S(n2206), .Y(n321) );
  INVX2 U666 ( .A(n321), .Y(n1844) );
  MUX2X1 U667 ( .B(core_block[760]), .A(n2152), .S(n2206), .Y(n322) );
  INVX2 U668 ( .A(n322), .Y(n1843) );
  MUX2X1 U669 ( .B(core_block[759]), .A(n2150), .S(n2206), .Y(n323) );
  INVX2 U670 ( .A(n323), .Y(n1842) );
  MUX2X1 U671 ( .B(core_block[758]), .A(n2148), .S(n2206), .Y(n324) );
  INVX2 U672 ( .A(n324), .Y(n1841) );
  MUX2X1 U673 ( .B(core_block[757]), .A(n2146), .S(n2206), .Y(n325) );
  INVX2 U674 ( .A(n325), .Y(n1840) );
  MUX2X1 U675 ( .B(core_block[756]), .A(n2144), .S(n2206), .Y(n326) );
  INVX2 U676 ( .A(n326), .Y(n1839) );
  MUX2X1 U677 ( .B(core_block[755]), .A(n2142), .S(n2206), .Y(n327) );
  INVX2 U678 ( .A(n327), .Y(n1838) );
  MUX2X1 U679 ( .B(core_block[754]), .A(n2140), .S(n2206), .Y(n328) );
  INVX2 U680 ( .A(n328), .Y(n1837) );
  MUX2X1 U681 ( .B(core_block[753]), .A(n2138), .S(n2206), .Y(n329) );
  INVX2 U682 ( .A(n329), .Y(n1836) );
  MUX2X1 U683 ( .B(core_block[752]), .A(n2136), .S(n2206), .Y(n330) );
  INVX2 U684 ( .A(n330), .Y(n1835) );
  MUX2X1 U685 ( .B(core_block[751]), .A(n2134), .S(n2206), .Y(n331) );
  INVX2 U686 ( .A(n331), .Y(n1834) );
  MUX2X1 U687 ( .B(core_block[750]), .A(n2132), .S(n2206), .Y(n332) );
  INVX2 U688 ( .A(n332), .Y(n1833) );
  MUX2X1 U689 ( .B(core_block[749]), .A(n2130), .S(n2206), .Y(n333) );
  INVX2 U690 ( .A(n333), .Y(n1832) );
  MUX2X1 U691 ( .B(core_block[748]), .A(n2128), .S(n2206), .Y(n334) );
  INVX2 U692 ( .A(n334), .Y(n1831) );
  MUX2X1 U693 ( .B(core_block[747]), .A(n2126), .S(n2206), .Y(n335) );
  INVX2 U694 ( .A(n335), .Y(n1830) );
  MUX2X1 U695 ( .B(core_block[746]), .A(n2124), .S(n2206), .Y(n336) );
  INVX2 U696 ( .A(n336), .Y(n1829) );
  MUX2X1 U697 ( .B(core_block[745]), .A(n2122), .S(n2206), .Y(n337) );
  INVX2 U698 ( .A(n337), .Y(n1828) );
  MUX2X1 U699 ( .B(core_block[744]), .A(n2120), .S(n2206), .Y(n338) );
  INVX2 U700 ( .A(n338), .Y(n1827) );
  MUX2X1 U701 ( .B(core_block[743]), .A(n2118), .S(n2206), .Y(n339) );
  INVX2 U702 ( .A(n339), .Y(n1826) );
  MUX2X1 U703 ( .B(core_block[742]), .A(n2116), .S(n2206), .Y(n340) );
  INVX2 U704 ( .A(n340), .Y(n1825) );
  MUX2X1 U705 ( .B(core_block[741]), .A(n2114), .S(n2206), .Y(n341) );
  INVX2 U706 ( .A(n341), .Y(n1824) );
  MUX2X1 U707 ( .B(core_block[740]), .A(n2112), .S(n2206), .Y(n342) );
  INVX2 U708 ( .A(n342), .Y(n1823) );
  MUX2X1 U709 ( .B(core_block[739]), .A(n2110), .S(n2206), .Y(n343) );
  INVX2 U710 ( .A(n343), .Y(n1822) );
  MUX2X1 U711 ( .B(core_block[738]), .A(n2108), .S(n2206), .Y(n344) );
  INVX2 U712 ( .A(n344), .Y(n1821) );
  MUX2X1 U713 ( .B(core_block[737]), .A(n2172), .S(n2206), .Y(n345) );
  INVX2 U714 ( .A(n345), .Y(n1820) );
  MUX2X1 U715 ( .B(core_block[736]), .A(n2170), .S(n2206), .Y(n346) );
  INVX2 U716 ( .A(n346), .Y(n1819) );
  MUX2X1 U717 ( .B(core_block[735]), .A(n2166), .S(n2204), .Y(n347) );
  INVX2 U718 ( .A(n347), .Y(n1818) );
  MUX2X1 U719 ( .B(core_block[734]), .A(n2164), .S(n2204), .Y(n348) );
  INVX2 U720 ( .A(n348), .Y(n1817) );
  MUX2X1 U721 ( .B(core_block[733]), .A(n2162), .S(n2204), .Y(n349) );
  INVX2 U722 ( .A(n349), .Y(n1816) );
  MUX2X1 U723 ( .B(core_block[732]), .A(n2160), .S(n2204), .Y(n350) );
  INVX2 U724 ( .A(n350), .Y(n1815) );
  MUX2X1 U725 ( .B(core_block[731]), .A(n2158), .S(n2204), .Y(n351) );
  INVX2 U726 ( .A(n351), .Y(n1814) );
  MUX2X1 U727 ( .B(core_block[730]), .A(n2156), .S(n2204), .Y(n352) );
  INVX2 U728 ( .A(n352), .Y(n1813) );
  MUX2X1 U729 ( .B(core_block[729]), .A(n2154), .S(n2204), .Y(n353) );
  INVX2 U730 ( .A(n353), .Y(n1812) );
  MUX2X1 U731 ( .B(core_block[728]), .A(n2152), .S(n2204), .Y(n354) );
  INVX2 U732 ( .A(n354), .Y(n1811) );
  MUX2X1 U733 ( .B(core_block[727]), .A(n2150), .S(n2204), .Y(n355) );
  INVX2 U734 ( .A(n355), .Y(n1810) );
  MUX2X1 U735 ( .B(core_block[726]), .A(n2148), .S(n2204), .Y(n356) );
  INVX2 U736 ( .A(n356), .Y(n1809) );
  MUX2X1 U737 ( .B(core_block[725]), .A(n2146), .S(n2204), .Y(n357) );
  INVX2 U738 ( .A(n357), .Y(n1808) );
  MUX2X1 U739 ( .B(core_block[724]), .A(n2144), .S(n2204), .Y(n358) );
  INVX2 U740 ( .A(n358), .Y(n1807) );
  MUX2X1 U741 ( .B(core_block[723]), .A(n2142), .S(n2204), .Y(n359) );
  INVX2 U742 ( .A(n359), .Y(n1806) );
  MUX2X1 U743 ( .B(core_block[722]), .A(n2140), .S(n2204), .Y(n360) );
  INVX2 U744 ( .A(n360), .Y(n1805) );
  MUX2X1 U745 ( .B(core_block[721]), .A(n2138), .S(n2204), .Y(n361) );
  INVX2 U746 ( .A(n361), .Y(n1804) );
  MUX2X1 U747 ( .B(core_block[720]), .A(n2136), .S(n2204), .Y(n362) );
  INVX2 U748 ( .A(n362), .Y(n1803) );
  MUX2X1 U749 ( .B(core_block[719]), .A(n2134), .S(n2204), .Y(n363) );
  INVX2 U750 ( .A(n363), .Y(n1802) );
  MUX2X1 U751 ( .B(core_block[718]), .A(n2132), .S(n2204), .Y(n364) );
  INVX2 U752 ( .A(n364), .Y(n1801) );
  MUX2X1 U753 ( .B(core_block[717]), .A(n2130), .S(n2204), .Y(n365) );
  INVX2 U754 ( .A(n365), .Y(n1800) );
  MUX2X1 U755 ( .B(core_block[716]), .A(n2128), .S(n2204), .Y(n366) );
  INVX2 U756 ( .A(n366), .Y(n1799) );
  MUX2X1 U757 ( .B(core_block[715]), .A(n2126), .S(n2204), .Y(n367) );
  INVX2 U758 ( .A(n367), .Y(n1798) );
  MUX2X1 U759 ( .B(core_block[714]), .A(n2124), .S(n2204), .Y(n368) );
  INVX2 U760 ( .A(n368), .Y(n1797) );
  MUX2X1 U761 ( .B(core_block[713]), .A(n2122), .S(n2204), .Y(n369) );
  INVX2 U762 ( .A(n369), .Y(n1796) );
  MUX2X1 U763 ( .B(core_block[712]), .A(n2120), .S(n2204), .Y(n370) );
  INVX2 U764 ( .A(n370), .Y(n1795) );
  MUX2X1 U765 ( .B(core_block[711]), .A(n2118), .S(n2204), .Y(n371) );
  INVX2 U766 ( .A(n371), .Y(n1794) );
  MUX2X1 U767 ( .B(core_block[710]), .A(n2116), .S(n2204), .Y(n372) );
  INVX2 U768 ( .A(n372), .Y(n1793) );
  MUX2X1 U769 ( .B(core_block[709]), .A(n2114), .S(n2204), .Y(n373) );
  INVX2 U770 ( .A(n373), .Y(n1792) );
  MUX2X1 U771 ( .B(core_block[708]), .A(n2112), .S(n2204), .Y(n374) );
  INVX2 U772 ( .A(n374), .Y(n1791) );
  MUX2X1 U773 ( .B(core_block[707]), .A(n2110), .S(n2204), .Y(n375) );
  INVX2 U774 ( .A(n375), .Y(n1790) );
  MUX2X1 U775 ( .B(core_block[706]), .A(n2108), .S(n2204), .Y(n376) );
  INVX2 U776 ( .A(n376), .Y(n1789) );
  MUX2X1 U777 ( .B(core_block[705]), .A(n2172), .S(n2204), .Y(n377) );
  INVX2 U778 ( .A(n377), .Y(n1788) );
  MUX2X1 U779 ( .B(core_block[704]), .A(n2170), .S(n2204), .Y(n378) );
  INVX2 U780 ( .A(n378), .Y(n1787) );
  MUX2X1 U781 ( .B(core_block[703]), .A(n2166), .S(n2202), .Y(n379) );
  INVX2 U782 ( .A(n379), .Y(n1786) );
  MUX2X1 U783 ( .B(core_block[702]), .A(n2164), .S(n2202), .Y(n380) );
  INVX2 U784 ( .A(n380), .Y(n1785) );
  MUX2X1 U785 ( .B(core_block[701]), .A(n2162), .S(n2202), .Y(n381) );
  INVX2 U786 ( .A(n381), .Y(n1784) );
  MUX2X1 U787 ( .B(core_block[700]), .A(n2160), .S(n2202), .Y(n382) );
  INVX2 U788 ( .A(n382), .Y(n1783) );
  MUX2X1 U789 ( .B(core_block[699]), .A(n2158), .S(n2202), .Y(n383) );
  INVX2 U790 ( .A(n383), .Y(n1782) );
  MUX2X1 U791 ( .B(core_block[698]), .A(n2156), .S(n2202), .Y(n384) );
  INVX2 U792 ( .A(n384), .Y(n1781) );
  MUX2X1 U793 ( .B(core_block[697]), .A(n2154), .S(n2202), .Y(n385) );
  INVX2 U794 ( .A(n385), .Y(n1780) );
  MUX2X1 U795 ( .B(core_block[696]), .A(n2152), .S(n2202), .Y(n386) );
  INVX2 U796 ( .A(n386), .Y(n1779) );
  MUX2X1 U797 ( .B(core_block[695]), .A(n2150), .S(n2202), .Y(n387) );
  INVX2 U798 ( .A(n387), .Y(n1778) );
  MUX2X1 U799 ( .B(core_block[694]), .A(n2148), .S(n2202), .Y(n388) );
  INVX2 U800 ( .A(n388), .Y(n1777) );
  MUX2X1 U801 ( .B(core_block[693]), .A(n2146), .S(n2202), .Y(n389) );
  INVX2 U802 ( .A(n389), .Y(n1776) );
  MUX2X1 U803 ( .B(core_block[692]), .A(n2144), .S(n2202), .Y(n390) );
  INVX2 U804 ( .A(n390), .Y(n1775) );
  MUX2X1 U805 ( .B(core_block[691]), .A(n2142), .S(n2202), .Y(n391) );
  INVX2 U806 ( .A(n391), .Y(n1774) );
  MUX2X1 U807 ( .B(core_block[690]), .A(n2140), .S(n2202), .Y(n392) );
  INVX2 U808 ( .A(n392), .Y(n1773) );
  MUX2X1 U809 ( .B(core_block[689]), .A(n2138), .S(n2202), .Y(n393) );
  INVX2 U810 ( .A(n393), .Y(n1772) );
  MUX2X1 U811 ( .B(core_block[688]), .A(n2136), .S(n2202), .Y(n394) );
  INVX2 U812 ( .A(n394), .Y(n1771) );
  MUX2X1 U813 ( .B(core_block[687]), .A(n2134), .S(n2202), .Y(n395) );
  INVX2 U814 ( .A(n395), .Y(n1770) );
  MUX2X1 U815 ( .B(core_block[686]), .A(n2132), .S(n2202), .Y(n396) );
  INVX2 U816 ( .A(n396), .Y(n1769) );
  MUX2X1 U817 ( .B(core_block[685]), .A(n2130), .S(n2202), .Y(n397) );
  INVX2 U818 ( .A(n397), .Y(n1768) );
  MUX2X1 U819 ( .B(core_block[684]), .A(n2128), .S(n2202), .Y(n398) );
  INVX2 U820 ( .A(n398), .Y(n1767) );
  MUX2X1 U821 ( .B(core_block[683]), .A(n2126), .S(n2202), .Y(n399) );
  INVX2 U822 ( .A(n399), .Y(n1766) );
  MUX2X1 U823 ( .B(core_block[682]), .A(n2124), .S(n2202), .Y(n400) );
  INVX2 U824 ( .A(n400), .Y(n1765) );
  MUX2X1 U825 ( .B(core_block[681]), .A(n2122), .S(n2202), .Y(n401) );
  INVX2 U826 ( .A(n401), .Y(n1764) );
  MUX2X1 U827 ( .B(core_block[680]), .A(n2120), .S(n2202), .Y(n402) );
  INVX2 U828 ( .A(n402), .Y(n1763) );
  MUX2X1 U829 ( .B(core_block[679]), .A(n2118), .S(n2202), .Y(n403) );
  INVX2 U830 ( .A(n403), .Y(n1762) );
  MUX2X1 U831 ( .B(core_block[678]), .A(n2116), .S(n2202), .Y(n404) );
  INVX2 U832 ( .A(n404), .Y(n1761) );
  MUX2X1 U833 ( .B(core_block[677]), .A(n2114), .S(n2202), .Y(n405) );
  INVX2 U834 ( .A(n405), .Y(n1760) );
  MUX2X1 U835 ( .B(core_block[676]), .A(n2112), .S(n2202), .Y(n406) );
  INVX2 U836 ( .A(n406), .Y(n1759) );
  MUX2X1 U837 ( .B(core_block[675]), .A(n2110), .S(n2202), .Y(n407) );
  INVX2 U838 ( .A(n407), .Y(n1758) );
  MUX2X1 U839 ( .B(core_block[674]), .A(n2108), .S(n2202), .Y(n408) );
  INVX2 U840 ( .A(n408), .Y(n1757) );
  MUX2X1 U841 ( .B(core_block[673]), .A(n2172), .S(n2202), .Y(n409) );
  INVX2 U842 ( .A(n409), .Y(n1756) );
  MUX2X1 U843 ( .B(core_block[672]), .A(n2170), .S(n2202), .Y(n410) );
  INVX2 U844 ( .A(n410), .Y(n1755) );
  MUX2X1 U845 ( .B(core_block[671]), .A(n2166), .S(n2200), .Y(n411) );
  INVX2 U846 ( .A(n411), .Y(n1754) );
  MUX2X1 U847 ( .B(core_block[670]), .A(n2164), .S(n2200), .Y(n412) );
  INVX2 U848 ( .A(n412), .Y(n1753) );
  MUX2X1 U849 ( .B(core_block[669]), .A(n2162), .S(n2200), .Y(n413) );
  INVX2 U850 ( .A(n413), .Y(n1752) );
  MUX2X1 U851 ( .B(core_block[668]), .A(n2160), .S(n2200), .Y(n414) );
  INVX2 U852 ( .A(n414), .Y(n1751) );
  MUX2X1 U853 ( .B(core_block[667]), .A(n2158), .S(n2200), .Y(n415) );
  INVX2 U854 ( .A(n415), .Y(n1750) );
  MUX2X1 U855 ( .B(core_block[666]), .A(n2156), .S(n2200), .Y(n416) );
  INVX2 U856 ( .A(n416), .Y(n1749) );
  MUX2X1 U857 ( .B(core_block[665]), .A(n2154), .S(n2200), .Y(n417) );
  INVX2 U858 ( .A(n417), .Y(n1748) );
  MUX2X1 U859 ( .B(core_block[664]), .A(n2152), .S(n2200), .Y(n418) );
  INVX2 U860 ( .A(n418), .Y(n1747) );
  MUX2X1 U861 ( .B(core_block[663]), .A(n2150), .S(n2200), .Y(n419) );
  INVX2 U862 ( .A(n419), .Y(n1746) );
  MUX2X1 U863 ( .B(core_block[662]), .A(n2148), .S(n2200), .Y(n420) );
  INVX2 U864 ( .A(n420), .Y(n1745) );
  MUX2X1 U865 ( .B(core_block[661]), .A(n2146), .S(n2200), .Y(n421) );
  INVX2 U866 ( .A(n421), .Y(n1744) );
  MUX2X1 U867 ( .B(core_block[660]), .A(n2144), .S(n2200), .Y(n422) );
  INVX2 U868 ( .A(n422), .Y(n1743) );
  MUX2X1 U869 ( .B(core_block[659]), .A(n2142), .S(n2200), .Y(n423) );
  INVX2 U870 ( .A(n423), .Y(n1742) );
  MUX2X1 U871 ( .B(core_block[658]), .A(n2140), .S(n2200), .Y(n424) );
  INVX2 U872 ( .A(n424), .Y(n1741) );
  MUX2X1 U873 ( .B(core_block[657]), .A(n2138), .S(n2200), .Y(n425) );
  INVX2 U874 ( .A(n425), .Y(n1740) );
  MUX2X1 U875 ( .B(core_block[656]), .A(n2136), .S(n2200), .Y(n426) );
  INVX2 U876 ( .A(n426), .Y(n1739) );
  MUX2X1 U877 ( .B(core_block[655]), .A(n2134), .S(n2200), .Y(n427) );
  INVX2 U878 ( .A(n427), .Y(n1738) );
  MUX2X1 U879 ( .B(core_block[654]), .A(n2132), .S(n2200), .Y(n428) );
  INVX2 U880 ( .A(n428), .Y(n1737) );
  MUX2X1 U881 ( .B(core_block[653]), .A(n2130), .S(n2200), .Y(n429) );
  INVX2 U882 ( .A(n429), .Y(n1736) );
  MUX2X1 U883 ( .B(core_block[652]), .A(n2128), .S(n2200), .Y(n430) );
  INVX2 U884 ( .A(n430), .Y(n1735) );
  MUX2X1 U885 ( .B(core_block[651]), .A(n2126), .S(n2200), .Y(n431) );
  INVX2 U886 ( .A(n431), .Y(n1734) );
  MUX2X1 U887 ( .B(core_block[650]), .A(n2124), .S(n2200), .Y(n432) );
  INVX2 U888 ( .A(n432), .Y(n1733) );
  MUX2X1 U889 ( .B(core_block[649]), .A(n2122), .S(n2200), .Y(n433) );
  INVX2 U890 ( .A(n433), .Y(n1732) );
  MUX2X1 U891 ( .B(core_block[648]), .A(n2120), .S(n2200), .Y(n434) );
  INVX2 U892 ( .A(n434), .Y(n1731) );
  MUX2X1 U893 ( .B(core_block[647]), .A(n2118), .S(n2200), .Y(n435) );
  INVX2 U894 ( .A(n435), .Y(n1730) );
  MUX2X1 U895 ( .B(core_block[646]), .A(n2116), .S(n2200), .Y(n436) );
  INVX2 U896 ( .A(n436), .Y(n1729) );
  MUX2X1 U897 ( .B(core_block[645]), .A(n2114), .S(n2200), .Y(n437) );
  INVX2 U898 ( .A(n437), .Y(n1728) );
  MUX2X1 U899 ( .B(core_block[644]), .A(n2112), .S(n2200), .Y(n438) );
  INVX2 U900 ( .A(n438), .Y(n1727) );
  MUX2X1 U901 ( .B(core_block[643]), .A(n2110), .S(n2200), .Y(n439) );
  INVX2 U902 ( .A(n439), .Y(n1726) );
  MUX2X1 U903 ( .B(core_block[642]), .A(n2108), .S(n2200), .Y(n440) );
  INVX2 U904 ( .A(n440), .Y(n1725) );
  MUX2X1 U905 ( .B(core_block[641]), .A(n2172), .S(n2200), .Y(n441) );
  INVX2 U906 ( .A(n441), .Y(n1724) );
  MUX2X1 U907 ( .B(core_block[640]), .A(n2170), .S(n2200), .Y(n442) );
  INVX2 U908 ( .A(n442), .Y(n1723) );
  MUX2X1 U909 ( .B(core_block[639]), .A(n2166), .S(n2198), .Y(n443) );
  INVX2 U910 ( .A(n443), .Y(n1722) );
  MUX2X1 U911 ( .B(core_block[638]), .A(n2164), .S(n2198), .Y(n444) );
  INVX2 U912 ( .A(n444), .Y(n1721) );
  MUX2X1 U913 ( .B(core_block[637]), .A(n2162), .S(n2198), .Y(n445) );
  INVX2 U914 ( .A(n445), .Y(n1720) );
  MUX2X1 U915 ( .B(core_block[636]), .A(n2160), .S(n2198), .Y(n446) );
  INVX2 U916 ( .A(n446), .Y(n1719) );
  MUX2X1 U917 ( .B(core_block[635]), .A(n2158), .S(n2198), .Y(n447) );
  INVX2 U918 ( .A(n447), .Y(n1718) );
  MUX2X1 U919 ( .B(core_block[634]), .A(n2156), .S(n2198), .Y(n448) );
  INVX2 U920 ( .A(n448), .Y(n1717) );
  MUX2X1 U921 ( .B(core_block[633]), .A(n2154), .S(n2198), .Y(n449) );
  INVX2 U922 ( .A(n449), .Y(n1716) );
  MUX2X1 U923 ( .B(core_block[632]), .A(n2152), .S(n2198), .Y(n450) );
  INVX2 U924 ( .A(n450), .Y(n1715) );
  MUX2X1 U925 ( .B(core_block[631]), .A(n2150), .S(n2198), .Y(n451) );
  INVX2 U926 ( .A(n451), .Y(n1714) );
  MUX2X1 U927 ( .B(core_block[630]), .A(n2148), .S(n2198), .Y(n452) );
  INVX2 U928 ( .A(n452), .Y(n1713) );
  MUX2X1 U929 ( .B(core_block[629]), .A(n2146), .S(n2198), .Y(n453) );
  INVX2 U930 ( .A(n453), .Y(n1712) );
  MUX2X1 U931 ( .B(core_block[628]), .A(n2144), .S(n2198), .Y(n454) );
  INVX2 U932 ( .A(n454), .Y(n1711) );
  MUX2X1 U933 ( .B(core_block[627]), .A(n2142), .S(n2198), .Y(n455) );
  INVX2 U934 ( .A(n455), .Y(n1710) );
  MUX2X1 U935 ( .B(core_block[626]), .A(n2140), .S(n2198), .Y(n456) );
  INVX2 U936 ( .A(n456), .Y(n1709) );
  MUX2X1 U937 ( .B(core_block[625]), .A(n2138), .S(n2198), .Y(n457) );
  INVX2 U938 ( .A(n457), .Y(n1708) );
  MUX2X1 U939 ( .B(core_block[624]), .A(n2136), .S(n2198), .Y(n458) );
  INVX2 U940 ( .A(n458), .Y(n1707) );
  MUX2X1 U941 ( .B(core_block[623]), .A(n2134), .S(n2198), .Y(n459) );
  INVX2 U942 ( .A(n459), .Y(n1706) );
  MUX2X1 U943 ( .B(core_block[622]), .A(n2132), .S(n2198), .Y(n460) );
  INVX2 U944 ( .A(n460), .Y(n1705) );
  MUX2X1 U945 ( .B(core_block[621]), .A(n2130), .S(n2198), .Y(n461) );
  INVX2 U946 ( .A(n461), .Y(n1704) );
  MUX2X1 U947 ( .B(core_block[620]), .A(n2128), .S(n2198), .Y(n462) );
  INVX2 U948 ( .A(n462), .Y(n1703) );
  MUX2X1 U949 ( .B(core_block[619]), .A(n2126), .S(n2198), .Y(n463) );
  INVX2 U950 ( .A(n463), .Y(n1702) );
  MUX2X1 U951 ( .B(core_block[618]), .A(n2124), .S(n2198), .Y(n464) );
  INVX2 U952 ( .A(n464), .Y(n1701) );
  MUX2X1 U953 ( .B(core_block[617]), .A(n2122), .S(n2198), .Y(n465) );
  INVX2 U954 ( .A(n465), .Y(n1700) );
  MUX2X1 U955 ( .B(core_block[616]), .A(n2120), .S(n2198), .Y(n466) );
  INVX2 U956 ( .A(n466), .Y(n1699) );
  MUX2X1 U957 ( .B(core_block[615]), .A(n2118), .S(n2198), .Y(n467) );
  INVX2 U958 ( .A(n467), .Y(n1698) );
  MUX2X1 U959 ( .B(core_block[614]), .A(n2116), .S(n2198), .Y(n468) );
  INVX2 U960 ( .A(n468), .Y(n1697) );
  MUX2X1 U961 ( .B(core_block[613]), .A(n2114), .S(n2198), .Y(n469) );
  INVX2 U962 ( .A(n469), .Y(n1696) );
  MUX2X1 U963 ( .B(core_block[612]), .A(n2112), .S(n2198), .Y(n470) );
  INVX2 U964 ( .A(n470), .Y(n1695) );
  MUX2X1 U965 ( .B(core_block[611]), .A(n2110), .S(n2198), .Y(n471) );
  INVX2 U966 ( .A(n471), .Y(n1694) );
  MUX2X1 U967 ( .B(core_block[610]), .A(n2108), .S(n2198), .Y(n472) );
  INVX2 U968 ( .A(n472), .Y(n1693) );
  MUX2X1 U969 ( .B(core_block[609]), .A(n2172), .S(n2198), .Y(n473) );
  INVX2 U970 ( .A(n473), .Y(n1692) );
  MUX2X1 U971 ( .B(core_block[608]), .A(n2170), .S(n2198), .Y(n474) );
  INVX2 U972 ( .A(n474), .Y(n1691) );
  MUX2X1 U973 ( .B(core_block[607]), .A(n2166), .S(n2196), .Y(n475) );
  INVX2 U974 ( .A(n475), .Y(n1690) );
  MUX2X1 U975 ( .B(core_block[606]), .A(n2164), .S(n2196), .Y(n476) );
  INVX2 U976 ( .A(n476), .Y(n1689) );
  MUX2X1 U977 ( .B(core_block[605]), .A(n2162), .S(n2196), .Y(n477) );
  INVX2 U978 ( .A(n477), .Y(n1688) );
  MUX2X1 U979 ( .B(core_block[604]), .A(n2160), .S(n2196), .Y(n478) );
  INVX2 U980 ( .A(n478), .Y(n1687) );
  MUX2X1 U981 ( .B(core_block[603]), .A(n2158), .S(n2196), .Y(n479) );
  INVX2 U982 ( .A(n479), .Y(n1686) );
  MUX2X1 U983 ( .B(core_block[602]), .A(n2156), .S(n2196), .Y(n480) );
  INVX2 U984 ( .A(n480), .Y(n1685) );
  MUX2X1 U985 ( .B(core_block[601]), .A(n2154), .S(n2196), .Y(n481) );
  INVX2 U986 ( .A(n481), .Y(n1684) );
  MUX2X1 U987 ( .B(core_block[600]), .A(n2152), .S(n2196), .Y(n482) );
  INVX2 U988 ( .A(n482), .Y(n1683) );
  MUX2X1 U989 ( .B(core_block[599]), .A(n2150), .S(n2196), .Y(n483) );
  INVX2 U990 ( .A(n483), .Y(n1682) );
  MUX2X1 U991 ( .B(core_block[598]), .A(n2148), .S(n2196), .Y(n484) );
  INVX2 U992 ( .A(n484), .Y(n1681) );
  MUX2X1 U993 ( .B(core_block[597]), .A(n2146), .S(n2196), .Y(n485) );
  INVX2 U994 ( .A(n485), .Y(n1680) );
  MUX2X1 U995 ( .B(core_block[596]), .A(n2144), .S(n2196), .Y(n486) );
  INVX2 U996 ( .A(n486), .Y(n1679) );
  MUX2X1 U997 ( .B(core_block[595]), .A(n2142), .S(n2196), .Y(n487) );
  INVX2 U998 ( .A(n487), .Y(n1678) );
  MUX2X1 U999 ( .B(core_block[594]), .A(n2140), .S(n2196), .Y(n488) );
  INVX2 U1000 ( .A(n488), .Y(n1677) );
  MUX2X1 U1001 ( .B(core_block[593]), .A(n2138), .S(n2196), .Y(n489) );
  INVX2 U1002 ( .A(n489), .Y(n1676) );
  MUX2X1 U1003 ( .B(core_block[592]), .A(n2136), .S(n2196), .Y(n490) );
  INVX2 U1004 ( .A(n490), .Y(n1675) );
  MUX2X1 U1005 ( .B(core_block[591]), .A(n2134), .S(n2196), .Y(n491) );
  INVX2 U1006 ( .A(n491), .Y(n1674) );
  MUX2X1 U1007 ( .B(core_block[590]), .A(n2132), .S(n2196), .Y(n492) );
  INVX2 U1008 ( .A(n492), .Y(n1673) );
  MUX2X1 U1009 ( .B(core_block[589]), .A(n2130), .S(n2196), .Y(n493) );
  INVX2 U1010 ( .A(n493), .Y(n1672) );
  MUX2X1 U1011 ( .B(core_block[588]), .A(n2128), .S(n2196), .Y(n494) );
  INVX2 U1012 ( .A(n494), .Y(n1671) );
  MUX2X1 U1013 ( .B(core_block[587]), .A(n2126), .S(n2196), .Y(n495) );
  INVX2 U1014 ( .A(n495), .Y(n1670) );
  MUX2X1 U1015 ( .B(core_block[586]), .A(n2124), .S(n2196), .Y(n496) );
  INVX2 U1016 ( .A(n496), .Y(n1669) );
  MUX2X1 U1017 ( .B(core_block[585]), .A(n2122), .S(n2196), .Y(n497) );
  INVX2 U1018 ( .A(n497), .Y(n1668) );
  MUX2X1 U1019 ( .B(core_block[584]), .A(n2120), .S(n2196), .Y(n498) );
  INVX2 U1020 ( .A(n498), .Y(n1667) );
  MUX2X1 U1021 ( .B(core_block[583]), .A(n2118), .S(n2196), .Y(n499) );
  INVX2 U1022 ( .A(n499), .Y(n1666) );
  MUX2X1 U1023 ( .B(core_block[582]), .A(n2116), .S(n2196), .Y(n500) );
  INVX2 U1024 ( .A(n500), .Y(n1665) );
  MUX2X1 U1025 ( .B(core_block[581]), .A(n2114), .S(n2196), .Y(n501) );
  INVX2 U1026 ( .A(n501), .Y(n1664) );
  MUX2X1 U1027 ( .B(core_block[580]), .A(n2112), .S(n2196), .Y(n502) );
  INVX2 U1028 ( .A(n502), .Y(n1663) );
  MUX2X1 U1029 ( .B(core_block[579]), .A(n2110), .S(n2196), .Y(n503) );
  INVX2 U1030 ( .A(n503), .Y(n1662) );
  MUX2X1 U1031 ( .B(core_block[578]), .A(n2108), .S(n2196), .Y(n504) );
  INVX2 U1032 ( .A(n504), .Y(n1661) );
  MUX2X1 U1033 ( .B(core_block[577]), .A(n2172), .S(n2196), .Y(n505) );
  INVX2 U1034 ( .A(n505), .Y(n1660) );
  MUX2X1 U1035 ( .B(core_block[576]), .A(n2170), .S(n2196), .Y(n506) );
  INVX2 U1036 ( .A(n506), .Y(n1659) );
  MUX2X1 U1037 ( .B(core_block[575]), .A(n2166), .S(n2194), .Y(n507) );
  INVX2 U1038 ( .A(n507), .Y(n1658) );
  MUX2X1 U1039 ( .B(core_block[574]), .A(n2164), .S(n2194), .Y(n508) );
  INVX2 U1040 ( .A(n508), .Y(n1657) );
  MUX2X1 U1041 ( .B(core_block[573]), .A(n2162), .S(n2194), .Y(n509) );
  INVX2 U1042 ( .A(n509), .Y(n1656) );
  MUX2X1 U1043 ( .B(core_block[572]), .A(n2160), .S(n2194), .Y(n510) );
  INVX2 U1044 ( .A(n510), .Y(n1655) );
  MUX2X1 U1045 ( .B(core_block[571]), .A(n2158), .S(n2194), .Y(n511) );
  INVX2 U1046 ( .A(n511), .Y(n1654) );
  MUX2X1 U1047 ( .B(core_block[570]), .A(n2156), .S(n2194), .Y(n512) );
  INVX2 U1048 ( .A(n512), .Y(n1653) );
  MUX2X1 U1049 ( .B(core_block[569]), .A(n2154), .S(n2194), .Y(n513) );
  INVX2 U1050 ( .A(n513), .Y(n1652) );
  MUX2X1 U1051 ( .B(core_block[568]), .A(n2152), .S(n2194), .Y(n514) );
  INVX2 U1052 ( .A(n514), .Y(n1651) );
  MUX2X1 U1053 ( .B(core_block[567]), .A(n2150), .S(n2194), .Y(n515) );
  INVX2 U1054 ( .A(n515), .Y(n1650) );
  MUX2X1 U1055 ( .B(core_block[566]), .A(n2148), .S(n2194), .Y(n516) );
  INVX2 U1056 ( .A(n516), .Y(n1649) );
  MUX2X1 U1057 ( .B(core_block[565]), .A(n2146), .S(n2194), .Y(n517) );
  INVX2 U1058 ( .A(n517), .Y(n1648) );
  MUX2X1 U1059 ( .B(core_block[564]), .A(n2144), .S(n2194), .Y(n518) );
  INVX2 U1060 ( .A(n518), .Y(n1647) );
  MUX2X1 U1061 ( .B(core_block[563]), .A(n2142), .S(n2194), .Y(n519) );
  INVX2 U1062 ( .A(n519), .Y(n1646) );
  MUX2X1 U1063 ( .B(core_block[562]), .A(n2140), .S(n2194), .Y(n520) );
  INVX2 U1064 ( .A(n520), .Y(n1645) );
  MUX2X1 U1065 ( .B(core_block[561]), .A(n2138), .S(n2194), .Y(n521) );
  INVX2 U1066 ( .A(n521), .Y(n1644) );
  MUX2X1 U1067 ( .B(core_block[560]), .A(n2136), .S(n2194), .Y(n522) );
  INVX2 U1068 ( .A(n522), .Y(n1643) );
  MUX2X1 U1069 ( .B(core_block[559]), .A(n2134), .S(n2194), .Y(n523) );
  INVX2 U1070 ( .A(n523), .Y(n1642) );
  MUX2X1 U1071 ( .B(core_block[558]), .A(n2132), .S(n2194), .Y(n524) );
  INVX2 U1072 ( .A(n524), .Y(n1641) );
  MUX2X1 U1073 ( .B(core_block[557]), .A(n2130), .S(n2194), .Y(n525) );
  INVX2 U1074 ( .A(n525), .Y(n1640) );
  MUX2X1 U1075 ( .B(core_block[556]), .A(n2128), .S(n2194), .Y(n526) );
  INVX2 U1076 ( .A(n526), .Y(n1639) );
  MUX2X1 U1077 ( .B(core_block[555]), .A(n2126), .S(n2194), .Y(n527) );
  INVX2 U1078 ( .A(n527), .Y(n1638) );
  MUX2X1 U1079 ( .B(core_block[554]), .A(n2124), .S(n2194), .Y(n528) );
  INVX2 U1080 ( .A(n528), .Y(n1637) );
  MUX2X1 U1081 ( .B(core_block[553]), .A(n2122), .S(n2194), .Y(n529) );
  INVX2 U1082 ( .A(n529), .Y(n1636) );
  MUX2X1 U1083 ( .B(core_block[552]), .A(n2120), .S(n2194), .Y(n530) );
  INVX2 U1084 ( .A(n530), .Y(n1635) );
  MUX2X1 U1085 ( .B(core_block[551]), .A(n2118), .S(n2194), .Y(n531) );
  INVX2 U1086 ( .A(n531), .Y(n1634) );
  MUX2X1 U1087 ( .B(core_block[550]), .A(n2116), .S(n2194), .Y(n532) );
  INVX2 U1088 ( .A(n532), .Y(n1633) );
  MUX2X1 U1089 ( .B(core_block[549]), .A(n2114), .S(n2194), .Y(n533) );
  INVX2 U1090 ( .A(n533), .Y(n1632) );
  MUX2X1 U1091 ( .B(core_block[548]), .A(n2112), .S(n2194), .Y(n534) );
  INVX2 U1092 ( .A(n534), .Y(n1631) );
  MUX2X1 U1093 ( .B(core_block[547]), .A(n2110), .S(n2194), .Y(n535) );
  INVX2 U1094 ( .A(n535), .Y(n1630) );
  MUX2X1 U1095 ( .B(core_block[546]), .A(n2108), .S(n2194), .Y(n536) );
  INVX2 U1096 ( .A(n536), .Y(n1629) );
  MUX2X1 U1097 ( .B(core_block[545]), .A(n2172), .S(n2194), .Y(n537) );
  INVX2 U1098 ( .A(n537), .Y(n1628) );
  MUX2X1 U1099 ( .B(core_block[544]), .A(n2170), .S(n2194), .Y(n538) );
  INVX2 U1100 ( .A(n538), .Y(n1627) );
  MUX2X1 U1101 ( .B(core_block[543]), .A(n2166), .S(n2192), .Y(n539) );
  INVX2 U1102 ( .A(n539), .Y(n1626) );
  MUX2X1 U1103 ( .B(core_block[542]), .A(n2164), .S(n2192), .Y(n540) );
  INVX2 U1104 ( .A(n540), .Y(n1625) );
  MUX2X1 U1105 ( .B(core_block[541]), .A(n2162), .S(n2192), .Y(n541) );
  INVX2 U1106 ( .A(n541), .Y(n1624) );
  MUX2X1 U1107 ( .B(core_block[540]), .A(n2160), .S(n2192), .Y(n542) );
  INVX2 U1108 ( .A(n542), .Y(n1623) );
  MUX2X1 U1109 ( .B(core_block[539]), .A(n2158), .S(n2192), .Y(n543) );
  INVX2 U1110 ( .A(n543), .Y(n1622) );
  MUX2X1 U1111 ( .B(core_block[538]), .A(n2156), .S(n2192), .Y(n544) );
  INVX2 U1112 ( .A(n544), .Y(n1621) );
  MUX2X1 U1113 ( .B(core_block[537]), .A(n2154), .S(n2192), .Y(n545) );
  INVX2 U1114 ( .A(n545), .Y(n1620) );
  MUX2X1 U1115 ( .B(core_block[536]), .A(n2152), .S(n2192), .Y(n546) );
  INVX2 U1116 ( .A(n546), .Y(n1619) );
  MUX2X1 U1117 ( .B(core_block[535]), .A(n2150), .S(n2192), .Y(n547) );
  INVX2 U1118 ( .A(n547), .Y(n1618) );
  MUX2X1 U1119 ( .B(core_block[534]), .A(n2148), .S(n2192), .Y(n548) );
  INVX2 U1120 ( .A(n548), .Y(n1617) );
  MUX2X1 U1121 ( .B(core_block[533]), .A(n2146), .S(n2192), .Y(n549) );
  INVX2 U1122 ( .A(n549), .Y(n1616) );
  MUX2X1 U1123 ( .B(core_block[532]), .A(n2144), .S(n2192), .Y(n550) );
  INVX2 U1124 ( .A(n550), .Y(n1615) );
  MUX2X1 U1125 ( .B(core_block[531]), .A(n2142), .S(n2192), .Y(n551) );
  INVX2 U1126 ( .A(n551), .Y(n1614) );
  MUX2X1 U1127 ( .B(core_block[530]), .A(n2140), .S(n2192), .Y(n552) );
  INVX2 U1128 ( .A(n552), .Y(n1613) );
  MUX2X1 U1129 ( .B(core_block[529]), .A(n2138), .S(n2192), .Y(n553) );
  INVX2 U1130 ( .A(n553), .Y(n1612) );
  MUX2X1 U1131 ( .B(core_block[528]), .A(n2136), .S(n2192), .Y(n554) );
  INVX2 U1132 ( .A(n554), .Y(n1611) );
  MUX2X1 U1133 ( .B(core_block[527]), .A(n2134), .S(n2192), .Y(n555) );
  INVX2 U1134 ( .A(n555), .Y(n1610) );
  MUX2X1 U1135 ( .B(core_block[526]), .A(n2132), .S(n2192), .Y(n556) );
  INVX2 U1136 ( .A(n556), .Y(n1609) );
  MUX2X1 U1137 ( .B(core_block[525]), .A(n2130), .S(n2192), .Y(n557) );
  INVX2 U1138 ( .A(n557), .Y(n1608) );
  MUX2X1 U1139 ( .B(core_block[524]), .A(n2128), .S(n2192), .Y(n558) );
  INVX2 U1140 ( .A(n558), .Y(n1607) );
  MUX2X1 U1141 ( .B(core_block[523]), .A(n2126), .S(n2192), .Y(n559) );
  INVX2 U1142 ( .A(n559), .Y(n1606) );
  MUX2X1 U1143 ( .B(core_block[522]), .A(n2124), .S(n2192), .Y(n560) );
  INVX2 U1144 ( .A(n560), .Y(n1605) );
  MUX2X1 U1145 ( .B(core_block[521]), .A(n2122), .S(n2192), .Y(n561) );
  INVX2 U1146 ( .A(n561), .Y(n1604) );
  MUX2X1 U1147 ( .B(core_block[520]), .A(n2120), .S(n2192), .Y(n562) );
  INVX2 U1148 ( .A(n562), .Y(n1603) );
  MUX2X1 U1149 ( .B(core_block[519]), .A(n2118), .S(n2192), .Y(n563) );
  INVX2 U1150 ( .A(n563), .Y(n1602) );
  MUX2X1 U1151 ( .B(core_block[518]), .A(n2116), .S(n2192), .Y(n564) );
  INVX2 U1152 ( .A(n564), .Y(n1601) );
  MUX2X1 U1153 ( .B(core_block[517]), .A(n2114), .S(n2192), .Y(n565) );
  INVX2 U1154 ( .A(n565), .Y(n1600) );
  MUX2X1 U1155 ( .B(core_block[516]), .A(n2112), .S(n2192), .Y(n566) );
  INVX2 U1156 ( .A(n566), .Y(n1599) );
  MUX2X1 U1157 ( .B(core_block[515]), .A(n2110), .S(n2192), .Y(n567) );
  INVX2 U1158 ( .A(n567), .Y(n1598) );
  MUX2X1 U1159 ( .B(core_block[514]), .A(n2108), .S(n2192), .Y(n568) );
  INVX2 U1160 ( .A(n568), .Y(n1597) );
  MUX2X1 U1161 ( .B(core_block[513]), .A(n2172), .S(n2192), .Y(n569) );
  INVX2 U1162 ( .A(n569), .Y(n1596) );
  MUX2X1 U1163 ( .B(core_block[512]), .A(n2170), .S(n2192), .Y(n570) );
  INVX2 U1164 ( .A(n570), .Y(n1595) );
  MUX2X1 U1165 ( .B(core_block[511]), .A(n2166), .S(n2190), .Y(n571) );
  INVX2 U1166 ( .A(n571), .Y(n1594) );
  MUX2X1 U1167 ( .B(core_block[510]), .A(n2164), .S(n2190), .Y(n572) );
  INVX2 U1168 ( .A(n572), .Y(n1593) );
  MUX2X1 U1169 ( .B(core_block[509]), .A(n2162), .S(n2190), .Y(n573) );
  INVX2 U1170 ( .A(n573), .Y(n1592) );
  MUX2X1 U1171 ( .B(core_block[508]), .A(n2160), .S(n2190), .Y(n574) );
  INVX2 U1172 ( .A(n574), .Y(n1591) );
  MUX2X1 U1173 ( .B(core_block[507]), .A(n2158), .S(n2190), .Y(n575) );
  INVX2 U1174 ( .A(n575), .Y(n1590) );
  MUX2X1 U1175 ( .B(core_block[506]), .A(n2156), .S(n2190), .Y(n576) );
  INVX2 U1176 ( .A(n576), .Y(n1589) );
  MUX2X1 U1177 ( .B(core_block[505]), .A(n2154), .S(n2190), .Y(n577) );
  INVX2 U1178 ( .A(n577), .Y(n1588) );
  MUX2X1 U1179 ( .B(core_block[504]), .A(n2152), .S(n2190), .Y(n578) );
  INVX2 U1180 ( .A(n578), .Y(n1587) );
  MUX2X1 U1181 ( .B(core_block[503]), .A(n2150), .S(n2190), .Y(n579) );
  INVX2 U1182 ( .A(n579), .Y(n1586) );
  MUX2X1 U1183 ( .B(core_block[502]), .A(n2148), .S(n2190), .Y(n580) );
  INVX2 U1184 ( .A(n580), .Y(n1585) );
  MUX2X1 U1185 ( .B(core_block[501]), .A(n2146), .S(n2190), .Y(n581) );
  INVX2 U1186 ( .A(n581), .Y(n1584) );
  MUX2X1 U1187 ( .B(core_block[500]), .A(n2144), .S(n2190), .Y(n582) );
  INVX2 U1188 ( .A(n582), .Y(n1583) );
  MUX2X1 U1189 ( .B(core_block[499]), .A(n2142), .S(n2190), .Y(n583) );
  INVX2 U1190 ( .A(n583), .Y(n1582) );
  MUX2X1 U1191 ( .B(core_block[498]), .A(n2140), .S(n2190), .Y(n584) );
  INVX2 U1192 ( .A(n584), .Y(n1581) );
  MUX2X1 U1193 ( .B(core_block[497]), .A(n2138), .S(n2190), .Y(n585) );
  INVX2 U1194 ( .A(n585), .Y(n1580) );
  MUX2X1 U1195 ( .B(core_block[496]), .A(n2136), .S(n2190), .Y(n586) );
  INVX2 U1196 ( .A(n586), .Y(n1579) );
  MUX2X1 U1197 ( .B(core_block[495]), .A(n2134), .S(n2190), .Y(n587) );
  INVX2 U1198 ( .A(n587), .Y(n1578) );
  MUX2X1 U1199 ( .B(core_block[494]), .A(n2132), .S(n2190), .Y(n588) );
  INVX2 U1200 ( .A(n588), .Y(n1577) );
  MUX2X1 U1201 ( .B(core_block[493]), .A(n2130), .S(n2190), .Y(n589) );
  INVX2 U1202 ( .A(n589), .Y(n1576) );
  MUX2X1 U1203 ( .B(core_block[492]), .A(n2128), .S(n2190), .Y(n590) );
  INVX2 U1204 ( .A(n590), .Y(n1575) );
  MUX2X1 U1205 ( .B(core_block[491]), .A(n2126), .S(n2190), .Y(n591) );
  INVX2 U1206 ( .A(n591), .Y(n1574) );
  MUX2X1 U1207 ( .B(core_block[490]), .A(n2124), .S(n2190), .Y(n592) );
  INVX2 U1208 ( .A(n592), .Y(n1573) );
  MUX2X1 U1209 ( .B(core_block[489]), .A(n2122), .S(n2190), .Y(n593) );
  INVX2 U1210 ( .A(n593), .Y(n1572) );
  MUX2X1 U1211 ( .B(core_block[488]), .A(n2120), .S(n2190), .Y(n594) );
  INVX2 U1212 ( .A(n594), .Y(n1571) );
  MUX2X1 U1213 ( .B(core_block[487]), .A(n2118), .S(n2190), .Y(n595) );
  INVX2 U1214 ( .A(n595), .Y(n1570) );
  MUX2X1 U1215 ( .B(core_block[486]), .A(n2116), .S(n2190), .Y(n596) );
  INVX2 U1216 ( .A(n596), .Y(n1569) );
  MUX2X1 U1217 ( .B(core_block[485]), .A(n2114), .S(n2190), .Y(n597) );
  INVX2 U1218 ( .A(n597), .Y(n1568) );
  MUX2X1 U1219 ( .B(core_block[484]), .A(n2112), .S(n2190), .Y(n598) );
  INVX2 U1220 ( .A(n598), .Y(n1567) );
  MUX2X1 U1221 ( .B(core_block[483]), .A(n2110), .S(n2190), .Y(n599) );
  INVX2 U1222 ( .A(n599), .Y(n1566) );
  MUX2X1 U1223 ( .B(core_block[482]), .A(n2108), .S(n2190), .Y(n600) );
  INVX2 U1224 ( .A(n600), .Y(n1565) );
  MUX2X1 U1225 ( .B(core_block[481]), .A(n2172), .S(n2190), .Y(n601) );
  INVX2 U1226 ( .A(n601), .Y(n1564) );
  MUX2X1 U1227 ( .B(core_block[480]), .A(n2170), .S(n2190), .Y(n602) );
  INVX2 U1228 ( .A(n602), .Y(n1563) );
  MUX2X1 U1229 ( .B(core_block[479]), .A(n2166), .S(n2188), .Y(n603) );
  INVX2 U1230 ( .A(n603), .Y(n1562) );
  MUX2X1 U1231 ( .B(core_block[478]), .A(n2164), .S(n2188), .Y(n604) );
  INVX2 U1232 ( .A(n604), .Y(n1561) );
  MUX2X1 U1233 ( .B(core_block[477]), .A(n2162), .S(n2188), .Y(n605) );
  INVX2 U1234 ( .A(n605), .Y(n1560) );
  MUX2X1 U1235 ( .B(core_block[476]), .A(n2160), .S(n2188), .Y(n606) );
  INVX2 U1236 ( .A(n606), .Y(n1559) );
  MUX2X1 U1237 ( .B(core_block[475]), .A(n2158), .S(n2188), .Y(n607) );
  INVX2 U1238 ( .A(n607), .Y(n1558) );
  MUX2X1 U1239 ( .B(core_block[474]), .A(n2156), .S(n2188), .Y(n608) );
  INVX2 U1240 ( .A(n608), .Y(n1557) );
  MUX2X1 U1241 ( .B(core_block[473]), .A(n2154), .S(n2188), .Y(n609) );
  INVX2 U1242 ( .A(n609), .Y(n1556) );
  MUX2X1 U1243 ( .B(core_block[472]), .A(n2152), .S(n2188), .Y(n610) );
  INVX2 U1244 ( .A(n610), .Y(n1555) );
  MUX2X1 U1245 ( .B(core_block[471]), .A(n2150), .S(n2188), .Y(n611) );
  INVX2 U1246 ( .A(n611), .Y(n1554) );
  MUX2X1 U1247 ( .B(core_block[470]), .A(n2148), .S(n2188), .Y(n612) );
  INVX2 U1248 ( .A(n612), .Y(n1553) );
  MUX2X1 U1249 ( .B(core_block[469]), .A(n2146), .S(n2188), .Y(n613) );
  INVX2 U1250 ( .A(n613), .Y(n1552) );
  MUX2X1 U1251 ( .B(core_block[468]), .A(n2144), .S(n2188), .Y(n614) );
  INVX2 U1252 ( .A(n614), .Y(n1551) );
  MUX2X1 U1253 ( .B(core_block[467]), .A(n2142), .S(n2188), .Y(n615) );
  INVX2 U1254 ( .A(n615), .Y(n1550) );
  MUX2X1 U1255 ( .B(core_block[466]), .A(n2140), .S(n2188), .Y(n616) );
  INVX2 U1256 ( .A(n616), .Y(n1549) );
  MUX2X1 U1257 ( .B(core_block[465]), .A(n2138), .S(n2188), .Y(n617) );
  INVX2 U1258 ( .A(n617), .Y(n1548) );
  MUX2X1 U1259 ( .B(core_block[464]), .A(n2136), .S(n2188), .Y(n618) );
  INVX2 U1260 ( .A(n618), .Y(n1547) );
  MUX2X1 U1261 ( .B(core_block[463]), .A(n2134), .S(n2188), .Y(n619) );
  INVX2 U1262 ( .A(n619), .Y(n1546) );
  MUX2X1 U1263 ( .B(core_block[462]), .A(n2132), .S(n2188), .Y(n620) );
  INVX2 U1264 ( .A(n620), .Y(n1545) );
  MUX2X1 U1265 ( .B(core_block[461]), .A(n2130), .S(n2188), .Y(n621) );
  INVX2 U1266 ( .A(n621), .Y(n1544) );
  MUX2X1 U1267 ( .B(core_block[460]), .A(n2128), .S(n2188), .Y(n622) );
  INVX2 U1268 ( .A(n622), .Y(n1543) );
  MUX2X1 U1269 ( .B(core_block[459]), .A(n2126), .S(n2188), .Y(n623) );
  INVX2 U1270 ( .A(n623), .Y(n1542) );
  MUX2X1 U1271 ( .B(core_block[458]), .A(n2124), .S(n2188), .Y(n624) );
  INVX2 U1272 ( .A(n624), .Y(n1541) );
  MUX2X1 U1273 ( .B(core_block[457]), .A(n2122), .S(n2188), .Y(n625) );
  INVX2 U1274 ( .A(n625), .Y(n1540) );
  MUX2X1 U1275 ( .B(core_block[456]), .A(n2120), .S(n2188), .Y(n626) );
  INVX2 U1276 ( .A(n626), .Y(n1539) );
  MUX2X1 U1277 ( .B(core_block[455]), .A(n2118), .S(n2188), .Y(n627) );
  INVX2 U1278 ( .A(n627), .Y(n1538) );
  MUX2X1 U1279 ( .B(core_block[454]), .A(n2116), .S(n2188), .Y(n628) );
  INVX2 U1280 ( .A(n628), .Y(n1537) );
  MUX2X1 U1281 ( .B(core_block[453]), .A(n2114), .S(n2188), .Y(n629) );
  INVX2 U1282 ( .A(n629), .Y(n1536) );
  MUX2X1 U1283 ( .B(core_block[452]), .A(n2112), .S(n2188), .Y(n630) );
  INVX2 U1284 ( .A(n630), .Y(n1535) );
  MUX2X1 U1285 ( .B(core_block[451]), .A(n2110), .S(n2188), .Y(n631) );
  INVX2 U1286 ( .A(n631), .Y(n1534) );
  MUX2X1 U1287 ( .B(core_block[450]), .A(n2108), .S(n2188), .Y(n632) );
  INVX2 U1288 ( .A(n632), .Y(n1533) );
  MUX2X1 U1289 ( .B(core_block[449]), .A(n2172), .S(n2188), .Y(n633) );
  INVX2 U1290 ( .A(n633), .Y(n1532) );
  MUX2X1 U1291 ( .B(core_block[448]), .A(n2170), .S(n2188), .Y(n634) );
  INVX2 U1292 ( .A(n634), .Y(n1531) );
  MUX2X1 U1293 ( .B(core_block[447]), .A(n2166), .S(n2186), .Y(n635) );
  INVX2 U1294 ( .A(n635), .Y(n1530) );
  MUX2X1 U1295 ( .B(core_block[446]), .A(n2164), .S(n2186), .Y(n636) );
  INVX2 U1296 ( .A(n636), .Y(n1529) );
  MUX2X1 U1297 ( .B(core_block[445]), .A(n2162), .S(n2186), .Y(n637) );
  INVX2 U1298 ( .A(n637), .Y(n1528) );
  MUX2X1 U1299 ( .B(core_block[444]), .A(n2160), .S(n2186), .Y(n638) );
  INVX2 U1300 ( .A(n638), .Y(n1527) );
  MUX2X1 U1301 ( .B(core_block[443]), .A(n2158), .S(n2186), .Y(n639) );
  INVX2 U1302 ( .A(n639), .Y(n1526) );
  MUX2X1 U1303 ( .B(core_block[442]), .A(n2156), .S(n2186), .Y(n640) );
  INVX2 U1304 ( .A(n640), .Y(n1525) );
  MUX2X1 U1305 ( .B(core_block[441]), .A(n2154), .S(n2186), .Y(n641) );
  INVX2 U1306 ( .A(n641), .Y(n1524) );
  MUX2X1 U1307 ( .B(core_block[440]), .A(n2152), .S(n2186), .Y(n642) );
  INVX2 U1308 ( .A(n642), .Y(n1523) );
  MUX2X1 U1309 ( .B(core_block[439]), .A(n2150), .S(n2186), .Y(n643) );
  INVX2 U1310 ( .A(n643), .Y(n1522) );
  MUX2X1 U1311 ( .B(core_block[438]), .A(n2148), .S(n2186), .Y(n644) );
  INVX2 U1312 ( .A(n644), .Y(n1521) );
  MUX2X1 U1313 ( .B(core_block[437]), .A(n2146), .S(n2186), .Y(n645) );
  INVX2 U1314 ( .A(n645), .Y(n1520) );
  MUX2X1 U1315 ( .B(core_block[436]), .A(n2144), .S(n2186), .Y(n646) );
  INVX2 U1316 ( .A(n646), .Y(n1519) );
  MUX2X1 U1317 ( .B(core_block[435]), .A(n2142), .S(n2186), .Y(n647) );
  INVX2 U1318 ( .A(n647), .Y(n1518) );
  MUX2X1 U1319 ( .B(core_block[434]), .A(n2140), .S(n2186), .Y(n648) );
  INVX2 U1320 ( .A(n648), .Y(n1517) );
  MUX2X1 U1321 ( .B(core_block[433]), .A(n2138), .S(n2186), .Y(n649) );
  INVX2 U1322 ( .A(n649), .Y(n1516) );
  MUX2X1 U1323 ( .B(core_block[432]), .A(n2136), .S(n2186), .Y(n650) );
  INVX2 U1324 ( .A(n650), .Y(n1515) );
  MUX2X1 U1325 ( .B(core_block[431]), .A(n2134), .S(n2186), .Y(n651) );
  INVX2 U1326 ( .A(n651), .Y(n1514) );
  MUX2X1 U1327 ( .B(core_block[430]), .A(n2132), .S(n2186), .Y(n652) );
  INVX2 U1328 ( .A(n652), .Y(n1513) );
  MUX2X1 U1329 ( .B(core_block[429]), .A(n2130), .S(n2186), .Y(n653) );
  INVX2 U1330 ( .A(n653), .Y(n1512) );
  MUX2X1 U1331 ( .B(core_block[428]), .A(n2128), .S(n2186), .Y(n654) );
  INVX2 U1332 ( .A(n654), .Y(n1511) );
  MUX2X1 U1333 ( .B(core_block[427]), .A(n2126), .S(n2186), .Y(n655) );
  INVX2 U1334 ( .A(n655), .Y(n1510) );
  MUX2X1 U1335 ( .B(core_block[426]), .A(n2124), .S(n2186), .Y(n656) );
  INVX2 U1336 ( .A(n656), .Y(n1509) );
  MUX2X1 U1337 ( .B(core_block[425]), .A(n2122), .S(n2186), .Y(n657) );
  INVX2 U1338 ( .A(n657), .Y(n1508) );
  MUX2X1 U1339 ( .B(core_block[424]), .A(n2120), .S(n2186), .Y(n658) );
  INVX2 U1340 ( .A(n658), .Y(n1507) );
  MUX2X1 U1341 ( .B(core_block[423]), .A(n2118), .S(n2186), .Y(n659) );
  INVX2 U1342 ( .A(n659), .Y(n1506) );
  MUX2X1 U1343 ( .B(core_block[422]), .A(n2116), .S(n2186), .Y(n660) );
  INVX2 U1344 ( .A(n660), .Y(n1505) );
  MUX2X1 U1345 ( .B(core_block[421]), .A(n2114), .S(n2186), .Y(n661) );
  INVX2 U1346 ( .A(n661), .Y(n1504) );
  MUX2X1 U1347 ( .B(core_block[420]), .A(n2112), .S(n2186), .Y(n662) );
  INVX2 U1348 ( .A(n662), .Y(n1503) );
  MUX2X1 U1349 ( .B(core_block[419]), .A(n2110), .S(n2186), .Y(n663) );
  INVX2 U1350 ( .A(n663), .Y(n1502) );
  MUX2X1 U1351 ( .B(core_block[418]), .A(n2108), .S(n2186), .Y(n664) );
  INVX2 U1352 ( .A(n664), .Y(n1501) );
  MUX2X1 U1353 ( .B(core_block[417]), .A(n2172), .S(n2186), .Y(n665) );
  INVX2 U1354 ( .A(n665), .Y(n1500) );
  MUX2X1 U1355 ( .B(core_block[416]), .A(n2170), .S(n2186), .Y(n666) );
  INVX2 U1356 ( .A(n666), .Y(n1499) );
  MUX2X1 U1357 ( .B(core_block[415]), .A(n2166), .S(n2184), .Y(n667) );
  INVX2 U1358 ( .A(n667), .Y(n1498) );
  MUX2X1 U1359 ( .B(core_block[414]), .A(n2164), .S(n2184), .Y(n668) );
  INVX2 U1360 ( .A(n668), .Y(n1497) );
  MUX2X1 U1361 ( .B(core_block[413]), .A(n2162), .S(n2184), .Y(n669) );
  INVX2 U1362 ( .A(n669), .Y(n1496) );
  MUX2X1 U1363 ( .B(core_block[412]), .A(n2160), .S(n2184), .Y(n670) );
  INVX2 U1364 ( .A(n670), .Y(n1495) );
  MUX2X1 U1365 ( .B(core_block[411]), .A(n2158), .S(n2184), .Y(n671) );
  INVX2 U1366 ( .A(n671), .Y(n1494) );
  MUX2X1 U1367 ( .B(core_block[410]), .A(n2156), .S(n2184), .Y(n672) );
  INVX2 U1368 ( .A(n672), .Y(n1493) );
  MUX2X1 U1369 ( .B(core_block[409]), .A(n2154), .S(n2184), .Y(n673) );
  INVX2 U1370 ( .A(n673), .Y(n1492) );
  MUX2X1 U1371 ( .B(core_block[408]), .A(n2152), .S(n2184), .Y(n674) );
  INVX2 U1372 ( .A(n674), .Y(n1491) );
  MUX2X1 U1373 ( .B(core_block[407]), .A(n2150), .S(n2184), .Y(n675) );
  INVX2 U1374 ( .A(n675), .Y(n1490) );
  MUX2X1 U1375 ( .B(core_block[406]), .A(n2148), .S(n2184), .Y(n676) );
  INVX2 U1376 ( .A(n676), .Y(n1489) );
  MUX2X1 U1377 ( .B(core_block[405]), .A(n2146), .S(n2184), .Y(n677) );
  INVX2 U1378 ( .A(n677), .Y(n1488) );
  MUX2X1 U1379 ( .B(core_block[404]), .A(n2144), .S(n2184), .Y(n678) );
  INVX2 U1380 ( .A(n678), .Y(n1487) );
  MUX2X1 U1381 ( .B(core_block[403]), .A(n2142), .S(n2184), .Y(n679) );
  INVX2 U1382 ( .A(n679), .Y(n1486) );
  MUX2X1 U1383 ( .B(core_block[402]), .A(n2140), .S(n2184), .Y(n680) );
  INVX2 U1384 ( .A(n680), .Y(n1485) );
  MUX2X1 U1385 ( .B(core_block[401]), .A(n2138), .S(n2184), .Y(n681) );
  INVX2 U1386 ( .A(n681), .Y(n1484) );
  MUX2X1 U1387 ( .B(core_block[400]), .A(n2136), .S(n2184), .Y(n682) );
  INVX2 U1388 ( .A(n682), .Y(n1483) );
  MUX2X1 U1389 ( .B(core_block[399]), .A(n2134), .S(n2184), .Y(n683) );
  INVX2 U1390 ( .A(n683), .Y(n1482) );
  MUX2X1 U1391 ( .B(core_block[398]), .A(n2132), .S(n2184), .Y(n684) );
  INVX2 U1392 ( .A(n684), .Y(n1481) );
  MUX2X1 U1393 ( .B(core_block[397]), .A(n2130), .S(n2184), .Y(n685) );
  INVX2 U1394 ( .A(n685), .Y(n1480) );
  MUX2X1 U1395 ( .B(core_block[396]), .A(n2128), .S(n2184), .Y(n686) );
  INVX2 U1396 ( .A(n686), .Y(n1479) );
  MUX2X1 U1397 ( .B(core_block[395]), .A(n2126), .S(n2184), .Y(n687) );
  INVX2 U1398 ( .A(n687), .Y(n1478) );
  MUX2X1 U1399 ( .B(core_block[394]), .A(n2124), .S(n2184), .Y(n688) );
  INVX2 U1400 ( .A(n688), .Y(n1477) );
  MUX2X1 U1401 ( .B(core_block[393]), .A(n2122), .S(n2184), .Y(n689) );
  INVX2 U1402 ( .A(n689), .Y(n1476) );
  MUX2X1 U1403 ( .B(core_block[392]), .A(n2120), .S(n2184), .Y(n690) );
  INVX2 U1404 ( .A(n690), .Y(n1475) );
  MUX2X1 U1405 ( .B(core_block[391]), .A(n2118), .S(n2184), .Y(n691) );
  INVX2 U1406 ( .A(n691), .Y(n1474) );
  MUX2X1 U1407 ( .B(core_block[390]), .A(n2116), .S(n2184), .Y(n692) );
  INVX2 U1408 ( .A(n692), .Y(n1473) );
  MUX2X1 U1409 ( .B(core_block[389]), .A(n2114), .S(n2184), .Y(n693) );
  INVX2 U1410 ( .A(n693), .Y(n1472) );
  MUX2X1 U1411 ( .B(core_block[388]), .A(n2112), .S(n2184), .Y(n694) );
  INVX2 U1412 ( .A(n694), .Y(n1471) );
  MUX2X1 U1413 ( .B(core_block[387]), .A(n2110), .S(n2184), .Y(n695) );
  INVX2 U1414 ( .A(n695), .Y(n1470) );
  MUX2X1 U1415 ( .B(core_block[386]), .A(n2108), .S(n2184), .Y(n696) );
  INVX2 U1416 ( .A(n696), .Y(n1469) );
  MUX2X1 U1417 ( .B(core_block[385]), .A(n2172), .S(n2184), .Y(n697) );
  INVX2 U1418 ( .A(n697), .Y(n1468) );
  MUX2X1 U1419 ( .B(core_block[384]), .A(n2170), .S(n2184), .Y(n698) );
  INVX2 U1420 ( .A(n698), .Y(n1467) );
  MUX2X1 U1421 ( .B(core_block[383]), .A(n2166), .S(n2182), .Y(n699) );
  INVX2 U1422 ( .A(n699), .Y(n1466) );
  MUX2X1 U1423 ( .B(core_block[382]), .A(n2164), .S(n2182), .Y(n700) );
  INVX2 U1424 ( .A(n700), .Y(n1465) );
  MUX2X1 U1425 ( .B(core_block[381]), .A(n2162), .S(n2182), .Y(n701) );
  INVX2 U1426 ( .A(n701), .Y(n1464) );
  MUX2X1 U1427 ( .B(core_block[380]), .A(n2160), .S(n2182), .Y(n702) );
  INVX2 U1428 ( .A(n702), .Y(n1463) );
  MUX2X1 U1429 ( .B(core_block[379]), .A(n2158), .S(n2182), .Y(n703) );
  INVX2 U1430 ( .A(n703), .Y(n1462) );
  MUX2X1 U1431 ( .B(core_block[378]), .A(n2156), .S(n2182), .Y(n704) );
  INVX2 U1432 ( .A(n704), .Y(n1461) );
  MUX2X1 U1433 ( .B(core_block[377]), .A(n2154), .S(n2182), .Y(n705) );
  INVX2 U1434 ( .A(n705), .Y(n1460) );
  MUX2X1 U1435 ( .B(core_block[376]), .A(n2152), .S(n2182), .Y(n706) );
  INVX2 U1436 ( .A(n706), .Y(n1459) );
  MUX2X1 U1437 ( .B(core_block[375]), .A(n2150), .S(n2182), .Y(n707) );
  INVX2 U1438 ( .A(n707), .Y(n1458) );
  MUX2X1 U1439 ( .B(core_block[374]), .A(n2148), .S(n2182), .Y(n708) );
  INVX2 U1440 ( .A(n708), .Y(n1457) );
  MUX2X1 U1441 ( .B(core_block[373]), .A(n2146), .S(n2182), .Y(n709) );
  INVX2 U1442 ( .A(n709), .Y(n1456) );
  MUX2X1 U1443 ( .B(core_block[372]), .A(n2144), .S(n2182), .Y(n710) );
  INVX2 U1444 ( .A(n710), .Y(n1455) );
  MUX2X1 U1445 ( .B(core_block[371]), .A(n2142), .S(n2182), .Y(n711) );
  INVX2 U1446 ( .A(n711), .Y(n1454) );
  MUX2X1 U1447 ( .B(core_block[370]), .A(n2140), .S(n2182), .Y(n712) );
  INVX2 U1448 ( .A(n712), .Y(n1453) );
  MUX2X1 U1449 ( .B(core_block[369]), .A(n2138), .S(n2182), .Y(n713) );
  INVX2 U1450 ( .A(n713), .Y(n1452) );
  MUX2X1 U1451 ( .B(core_block[368]), .A(n2136), .S(n2182), .Y(n714) );
  INVX2 U1452 ( .A(n714), .Y(n1451) );
  MUX2X1 U1453 ( .B(core_block[367]), .A(n2134), .S(n2182), .Y(n715) );
  INVX2 U1454 ( .A(n715), .Y(n1450) );
  MUX2X1 U1455 ( .B(core_block[366]), .A(n2132), .S(n2182), .Y(n716) );
  INVX2 U1456 ( .A(n716), .Y(n1449) );
  MUX2X1 U1457 ( .B(core_block[365]), .A(n2130), .S(n2182), .Y(n717) );
  INVX2 U1458 ( .A(n717), .Y(n1448) );
  MUX2X1 U1459 ( .B(core_block[364]), .A(n2128), .S(n2182), .Y(n718) );
  INVX2 U1460 ( .A(n718), .Y(n1447) );
  MUX2X1 U1461 ( .B(core_block[363]), .A(n2126), .S(n2182), .Y(n719) );
  INVX2 U1462 ( .A(n719), .Y(n1446) );
  MUX2X1 U1463 ( .B(core_block[362]), .A(n2124), .S(n2182), .Y(n720) );
  INVX2 U1464 ( .A(n720), .Y(n1445) );
  MUX2X1 U1465 ( .B(core_block[361]), .A(n2122), .S(n2182), .Y(n721) );
  INVX2 U1466 ( .A(n721), .Y(n1444) );
  MUX2X1 U1467 ( .B(core_block[360]), .A(n2120), .S(n2182), .Y(n722) );
  INVX2 U1468 ( .A(n722), .Y(n1443) );
  MUX2X1 U1469 ( .B(core_block[359]), .A(n2118), .S(n2182), .Y(n723) );
  INVX2 U1470 ( .A(n723), .Y(n1442) );
  MUX2X1 U1471 ( .B(core_block[358]), .A(n2116), .S(n2182), .Y(n724) );
  INVX2 U1472 ( .A(n724), .Y(n1441) );
  MUX2X1 U1473 ( .B(core_block[357]), .A(n2114), .S(n2182), .Y(n725) );
  INVX2 U1474 ( .A(n725), .Y(n1440) );
  MUX2X1 U1475 ( .B(core_block[356]), .A(n2112), .S(n2182), .Y(n726) );
  INVX2 U1476 ( .A(n726), .Y(n1439) );
  MUX2X1 U1477 ( .B(core_block[355]), .A(n2110), .S(n2182), .Y(n727) );
  INVX2 U1478 ( .A(n727), .Y(n1438) );
  MUX2X1 U1479 ( .B(core_block[354]), .A(n2108), .S(n2182), .Y(n728) );
  INVX2 U1480 ( .A(n728), .Y(n1437) );
  MUX2X1 U1481 ( .B(core_block[353]), .A(n2172), .S(n2182), .Y(n729) );
  INVX2 U1482 ( .A(n729), .Y(n1436) );
  MUX2X1 U1483 ( .B(core_block[352]), .A(n2170), .S(n2182), .Y(n730) );
  INVX2 U1484 ( .A(n730), .Y(n1435) );
  MUX2X1 U1485 ( .B(core_block[351]), .A(n2166), .S(n2180), .Y(n731) );
  INVX2 U1486 ( .A(n731), .Y(n1434) );
  MUX2X1 U1487 ( .B(core_block[350]), .A(n2164), .S(n2180), .Y(n732) );
  INVX2 U1488 ( .A(n732), .Y(n1433) );
  MUX2X1 U1489 ( .B(core_block[349]), .A(n2162), .S(n2180), .Y(n733) );
  INVX2 U1490 ( .A(n733), .Y(n1432) );
  MUX2X1 U1491 ( .B(core_block[348]), .A(n2160), .S(n2180), .Y(n734) );
  INVX2 U1492 ( .A(n734), .Y(n1431) );
  MUX2X1 U1493 ( .B(core_block[347]), .A(n2158), .S(n2180), .Y(n735) );
  INVX2 U1494 ( .A(n735), .Y(n1430) );
  MUX2X1 U1495 ( .B(core_block[346]), .A(n2156), .S(n2180), .Y(n736) );
  INVX2 U1496 ( .A(n736), .Y(n1429) );
  MUX2X1 U1497 ( .B(core_block[345]), .A(n2154), .S(n2180), .Y(n737) );
  INVX2 U1498 ( .A(n737), .Y(n1428) );
  MUX2X1 U1499 ( .B(core_block[344]), .A(n2152), .S(n2180), .Y(n738) );
  INVX2 U1500 ( .A(n738), .Y(n1427) );
  MUX2X1 U1501 ( .B(core_block[343]), .A(n2150), .S(n2180), .Y(n739) );
  INVX2 U1502 ( .A(n739), .Y(n1426) );
  MUX2X1 U1503 ( .B(core_block[342]), .A(n2148), .S(n2180), .Y(n740) );
  INVX2 U1504 ( .A(n740), .Y(n1425) );
  MUX2X1 U1505 ( .B(core_block[341]), .A(n2146), .S(n2180), .Y(n741) );
  INVX2 U1506 ( .A(n741), .Y(n1424) );
  MUX2X1 U1507 ( .B(core_block[340]), .A(n2144), .S(n2180), .Y(n742) );
  INVX2 U1508 ( .A(n742), .Y(n1423) );
  MUX2X1 U1509 ( .B(core_block[339]), .A(n2142), .S(n2180), .Y(n743) );
  INVX2 U1510 ( .A(n743), .Y(n1422) );
  MUX2X1 U1511 ( .B(core_block[338]), .A(n2140), .S(n2180), .Y(n744) );
  INVX2 U1512 ( .A(n744), .Y(n1421) );
  MUX2X1 U1513 ( .B(core_block[337]), .A(n2138), .S(n2180), .Y(n745) );
  INVX2 U1514 ( .A(n745), .Y(n1420) );
  MUX2X1 U1515 ( .B(core_block[336]), .A(n2136), .S(n2180), .Y(n746) );
  INVX2 U1516 ( .A(n746), .Y(n1419) );
  MUX2X1 U1517 ( .B(core_block[335]), .A(n2134), .S(n2180), .Y(n747) );
  INVX2 U1518 ( .A(n747), .Y(n1418) );
  MUX2X1 U1519 ( .B(core_block[334]), .A(n2132), .S(n2180), .Y(n748) );
  INVX2 U1520 ( .A(n748), .Y(n1417) );
  MUX2X1 U1521 ( .B(core_block[333]), .A(n2130), .S(n2180), .Y(n749) );
  INVX2 U1522 ( .A(n749), .Y(n1416) );
  MUX2X1 U1523 ( .B(core_block[332]), .A(n2128), .S(n2180), .Y(n750) );
  INVX2 U1524 ( .A(n750), .Y(n1415) );
  MUX2X1 U1525 ( .B(core_block[331]), .A(n2126), .S(n2180), .Y(n751) );
  INVX2 U1526 ( .A(n751), .Y(n1414) );
  MUX2X1 U1527 ( .B(core_block[330]), .A(n2124), .S(n2180), .Y(n752) );
  INVX2 U1528 ( .A(n752), .Y(n1413) );
  MUX2X1 U1529 ( .B(core_block[329]), .A(n2122), .S(n2180), .Y(n753) );
  INVX2 U1530 ( .A(n753), .Y(n1412) );
  MUX2X1 U1531 ( .B(core_block[328]), .A(n2120), .S(n2180), .Y(n754) );
  INVX2 U1532 ( .A(n754), .Y(n1411) );
  MUX2X1 U1533 ( .B(core_block[327]), .A(n2118), .S(n2180), .Y(n755) );
  INVX2 U1534 ( .A(n755), .Y(n1410) );
  MUX2X1 U1535 ( .B(core_block[326]), .A(n2116), .S(n2180), .Y(n756) );
  INVX2 U1536 ( .A(n756), .Y(n1409) );
  MUX2X1 U1537 ( .B(core_block[325]), .A(n2114), .S(n2180), .Y(n757) );
  INVX2 U1538 ( .A(n757), .Y(n1408) );
  MUX2X1 U1539 ( .B(core_block[324]), .A(n2112), .S(n2180), .Y(n758) );
  INVX2 U1540 ( .A(n758), .Y(n1407) );
  MUX2X1 U1541 ( .B(core_block[323]), .A(n2110), .S(n2180), .Y(n759) );
  INVX2 U1542 ( .A(n759), .Y(n1406) );
  MUX2X1 U1543 ( .B(core_block[322]), .A(n2108), .S(n2180), .Y(n760) );
  INVX2 U1544 ( .A(n760), .Y(n1405) );
  MUX2X1 U1545 ( .B(core_block[321]), .A(n2172), .S(n2180), .Y(n761) );
  INVX2 U1546 ( .A(n761), .Y(n1404) );
  MUX2X1 U1547 ( .B(core_block[320]), .A(n2170), .S(n2180), .Y(n762) );
  INVX2 U1548 ( .A(n762), .Y(n1403) );
  MUX2X1 U1549 ( .B(core_block[319]), .A(n2166), .S(n2178), .Y(n763) );
  INVX2 U1550 ( .A(n763), .Y(n1402) );
  MUX2X1 U1551 ( .B(core_block[318]), .A(n2164), .S(n2178), .Y(n764) );
  INVX2 U1552 ( .A(n764), .Y(n1401) );
  MUX2X1 U1553 ( .B(core_block[317]), .A(n2162), .S(n2178), .Y(n765) );
  INVX2 U1554 ( .A(n765), .Y(n1400) );
  MUX2X1 U1555 ( .B(core_block[316]), .A(n2160), .S(n2178), .Y(n766) );
  INVX2 U1556 ( .A(n766), .Y(n1399) );
  MUX2X1 U1557 ( .B(core_block[315]), .A(n2158), .S(n2178), .Y(n767) );
  INVX2 U1558 ( .A(n767), .Y(n1398) );
  MUX2X1 U1559 ( .B(core_block[314]), .A(n2156), .S(n2178), .Y(n768) );
  INVX2 U1560 ( .A(n768), .Y(n1397) );
  MUX2X1 U1561 ( .B(core_block[313]), .A(n2154), .S(n2178), .Y(n769) );
  INVX2 U1562 ( .A(n769), .Y(n1396) );
  MUX2X1 U1563 ( .B(core_block[312]), .A(n2152), .S(n2178), .Y(n770) );
  INVX2 U1564 ( .A(n770), .Y(n1395) );
  MUX2X1 U1565 ( .B(core_block[311]), .A(n2150), .S(n2178), .Y(n771) );
  INVX2 U1566 ( .A(n771), .Y(n1394) );
  MUX2X1 U1567 ( .B(core_block[310]), .A(n2148), .S(n2178), .Y(n772) );
  INVX2 U1568 ( .A(n772), .Y(n1393) );
  MUX2X1 U1569 ( .B(core_block[309]), .A(n2146), .S(n2178), .Y(n773) );
  INVX2 U1570 ( .A(n773), .Y(n1392) );
  MUX2X1 U1571 ( .B(core_block[308]), .A(n2144), .S(n2178), .Y(n774) );
  INVX2 U1572 ( .A(n774), .Y(n1391) );
  MUX2X1 U1573 ( .B(core_block[307]), .A(n2142), .S(n2178), .Y(n775) );
  INVX2 U1574 ( .A(n775), .Y(n1390) );
  MUX2X1 U1575 ( .B(core_block[306]), .A(n2140), .S(n2178), .Y(n776) );
  INVX2 U1576 ( .A(n776), .Y(n1389) );
  MUX2X1 U1577 ( .B(core_block[305]), .A(n2138), .S(n2178), .Y(n777) );
  INVX2 U1578 ( .A(n777), .Y(n1388) );
  MUX2X1 U1579 ( .B(core_block[304]), .A(n2136), .S(n2178), .Y(n778) );
  INVX2 U1580 ( .A(n778), .Y(n1387) );
  MUX2X1 U1581 ( .B(core_block[303]), .A(n2134), .S(n2178), .Y(n779) );
  INVX2 U1582 ( .A(n779), .Y(n1386) );
  MUX2X1 U1583 ( .B(core_block[302]), .A(n2132), .S(n2178), .Y(n780) );
  INVX2 U1584 ( .A(n780), .Y(n1385) );
  MUX2X1 U1585 ( .B(core_block[301]), .A(n2130), .S(n2178), .Y(n781) );
  INVX2 U1586 ( .A(n781), .Y(n1384) );
  MUX2X1 U1587 ( .B(core_block[300]), .A(n2128), .S(n2178), .Y(n782) );
  INVX2 U1588 ( .A(n782), .Y(n1383) );
  MUX2X1 U1589 ( .B(core_block[299]), .A(n2126), .S(n2178), .Y(n783) );
  INVX2 U1590 ( .A(n783), .Y(n1382) );
  MUX2X1 U1591 ( .B(core_block[298]), .A(n2124), .S(n2178), .Y(n784) );
  INVX2 U1592 ( .A(n784), .Y(n1381) );
  MUX2X1 U1593 ( .B(core_block[297]), .A(n2122), .S(n2178), .Y(n785) );
  INVX2 U1594 ( .A(n785), .Y(n1380) );
  MUX2X1 U1595 ( .B(core_block[296]), .A(n2120), .S(n2178), .Y(n786) );
  INVX2 U1596 ( .A(n786), .Y(n1379) );
  MUX2X1 U1597 ( .B(core_block[295]), .A(n2118), .S(n2178), .Y(n787) );
  INVX2 U1598 ( .A(n787), .Y(n1378) );
  MUX2X1 U1599 ( .B(core_block[294]), .A(n2116), .S(n2178), .Y(n788) );
  INVX2 U1600 ( .A(n788), .Y(n1377) );
  MUX2X1 U1601 ( .B(core_block[293]), .A(n2114), .S(n2178), .Y(n789) );
  INVX2 U1602 ( .A(n789), .Y(n1376) );
  MUX2X1 U1603 ( .B(core_block[292]), .A(n2112), .S(n2178), .Y(n790) );
  INVX2 U1604 ( .A(n790), .Y(n1375) );
  MUX2X1 U1605 ( .B(core_block[291]), .A(n2110), .S(n2178), .Y(n791) );
  INVX2 U1606 ( .A(n791), .Y(n1374) );
  MUX2X1 U1607 ( .B(core_block[290]), .A(n2108), .S(n2178), .Y(n792) );
  INVX2 U1608 ( .A(n792), .Y(n1373) );
  MUX2X1 U1609 ( .B(core_block[289]), .A(n2172), .S(n2178), .Y(n793) );
  INVX2 U1610 ( .A(n793), .Y(n1372) );
  MUX2X1 U1611 ( .B(core_block[288]), .A(n2170), .S(n2178), .Y(n794) );
  INVX2 U1612 ( .A(n794), .Y(n1371) );
  MUX2X1 U1613 ( .B(core_block[287]), .A(n2166), .S(n2176), .Y(n795) );
  INVX2 U1614 ( .A(n795), .Y(n1370) );
  MUX2X1 U1615 ( .B(core_block[286]), .A(n2164), .S(n2176), .Y(n796) );
  INVX2 U1616 ( .A(n796), .Y(n1369) );
  MUX2X1 U1617 ( .B(core_block[285]), .A(n2162), .S(n2176), .Y(n797) );
  INVX2 U1618 ( .A(n797), .Y(n1368) );
  MUX2X1 U1619 ( .B(core_block[284]), .A(n2160), .S(n2176), .Y(n798) );
  INVX2 U1620 ( .A(n798), .Y(n1367) );
  MUX2X1 U1621 ( .B(core_block[283]), .A(n2158), .S(n2176), .Y(n799) );
  INVX2 U1622 ( .A(n799), .Y(n1366) );
  MUX2X1 U1623 ( .B(core_block[282]), .A(n2156), .S(n2176), .Y(n800) );
  INVX2 U1624 ( .A(n800), .Y(n1365) );
  MUX2X1 U1625 ( .B(core_block[281]), .A(n2154), .S(n2176), .Y(n801) );
  INVX2 U1626 ( .A(n801), .Y(n1364) );
  MUX2X1 U1627 ( .B(core_block[280]), .A(n2152), .S(n2176), .Y(n802) );
  INVX2 U1628 ( .A(n802), .Y(n1363) );
  MUX2X1 U1629 ( .B(core_block[279]), .A(n2150), .S(n2176), .Y(n803) );
  INVX2 U1630 ( .A(n803), .Y(n1362) );
  MUX2X1 U1631 ( .B(core_block[278]), .A(n2148), .S(n2176), .Y(n804) );
  INVX2 U1632 ( .A(n804), .Y(n1361) );
  MUX2X1 U1633 ( .B(core_block[277]), .A(n2146), .S(n2176), .Y(n805) );
  INVX2 U1634 ( .A(n805), .Y(n1360) );
  MUX2X1 U1635 ( .B(core_block[276]), .A(n2144), .S(n2176), .Y(n806) );
  INVX2 U1636 ( .A(n806), .Y(n1359) );
  MUX2X1 U1637 ( .B(core_block[275]), .A(n2142), .S(n2176), .Y(n807) );
  INVX2 U1638 ( .A(n807), .Y(n1358) );
  MUX2X1 U1639 ( .B(core_block[274]), .A(n2140), .S(n2176), .Y(n808) );
  INVX2 U1640 ( .A(n808), .Y(n1357) );
  MUX2X1 U1641 ( .B(core_block[273]), .A(n2138), .S(n2176), .Y(n809) );
  INVX2 U1642 ( .A(n809), .Y(n1356) );
  MUX2X1 U1643 ( .B(core_block[272]), .A(n2136), .S(n2176), .Y(n810) );
  INVX2 U1644 ( .A(n810), .Y(n1355) );
  MUX2X1 U1645 ( .B(core_block[271]), .A(n2134), .S(n2176), .Y(n811) );
  INVX2 U1646 ( .A(n811), .Y(n1354) );
  MUX2X1 U1647 ( .B(core_block[270]), .A(n2132), .S(n2176), .Y(n812) );
  INVX2 U1648 ( .A(n812), .Y(n1353) );
  MUX2X1 U1649 ( .B(core_block[269]), .A(n2130), .S(n2176), .Y(n813) );
  INVX2 U1650 ( .A(n813), .Y(n1352) );
  MUX2X1 U1651 ( .B(core_block[268]), .A(n2128), .S(n2176), .Y(n814) );
  INVX2 U1652 ( .A(n814), .Y(n1351) );
  MUX2X1 U1653 ( .B(core_block[267]), .A(n2126), .S(n2176), .Y(n815) );
  INVX2 U1654 ( .A(n815), .Y(n1350) );
  MUX2X1 U1655 ( .B(core_block[266]), .A(n2124), .S(n2176), .Y(n816) );
  INVX2 U1656 ( .A(n816), .Y(n1349) );
  MUX2X1 U1657 ( .B(core_block[265]), .A(n2122), .S(n2176), .Y(n817) );
  INVX2 U1658 ( .A(n817), .Y(n1348) );
  MUX2X1 U1659 ( .B(core_block[264]), .A(n2120), .S(n2176), .Y(n818) );
  INVX2 U1660 ( .A(n818), .Y(n1347) );
  MUX2X1 U1661 ( .B(core_block[263]), .A(n2118), .S(n2176), .Y(n819) );
  INVX2 U1662 ( .A(n819), .Y(n1346) );
  MUX2X1 U1663 ( .B(core_block[262]), .A(n2116), .S(n2176), .Y(n820) );
  INVX2 U1664 ( .A(n820), .Y(n1345) );
  MUX2X1 U1665 ( .B(core_block[261]), .A(n2114), .S(n2176), .Y(n821) );
  INVX2 U1666 ( .A(n821), .Y(n1344) );
  MUX2X1 U1667 ( .B(core_block[260]), .A(n2112), .S(n2176), .Y(n822) );
  INVX2 U1668 ( .A(n822), .Y(n1343) );
  MUX2X1 U1669 ( .B(core_block[259]), .A(n2110), .S(n2176), .Y(n823) );
  INVX2 U1670 ( .A(n823), .Y(n1342) );
  MUX2X1 U1671 ( .B(core_block[258]), .A(n2108), .S(n2176), .Y(n824) );
  INVX2 U1672 ( .A(n824), .Y(n1341) );
  MUX2X1 U1673 ( .B(core_block[257]), .A(n2172), .S(n2176), .Y(n825) );
  INVX2 U1674 ( .A(n825), .Y(n1340) );
  MUX2X1 U1675 ( .B(core_block[256]), .A(n2170), .S(n2176), .Y(n826) );
  INVX2 U1676 ( .A(n826), .Y(n1339) );
  MUX2X1 U1677 ( .B(core_block[255]), .A(n2166), .S(n2174), .Y(n827) );
  INVX2 U1678 ( .A(n827), .Y(n1338) );
  MUX2X1 U1679 ( .B(core_block[254]), .A(n2164), .S(n2174), .Y(n828) );
  INVX2 U1680 ( .A(n828), .Y(n1337) );
  MUX2X1 U1681 ( .B(core_block[253]), .A(n2162), .S(n2174), .Y(n829) );
  INVX2 U1682 ( .A(n829), .Y(n1336) );
  MUX2X1 U1683 ( .B(core_block[252]), .A(n2160), .S(n2174), .Y(n830) );
  INVX2 U1684 ( .A(n830), .Y(n1335) );
  MUX2X1 U1685 ( .B(core_block[251]), .A(n2158), .S(n2174), .Y(n831) );
  INVX2 U1686 ( .A(n831), .Y(n1334) );
  MUX2X1 U1687 ( .B(core_block[250]), .A(n2156), .S(n2174), .Y(n832) );
  INVX2 U1688 ( .A(n832), .Y(n1333) );
  MUX2X1 U1689 ( .B(core_block[249]), .A(n2154), .S(n2174), .Y(n833) );
  INVX2 U1690 ( .A(n833), .Y(n1332) );
  MUX2X1 U1691 ( .B(core_block[248]), .A(n2152), .S(n2174), .Y(n834) );
  INVX2 U1692 ( .A(n834), .Y(n1331) );
  MUX2X1 U1693 ( .B(core_block[247]), .A(n2150), .S(n2174), .Y(n835) );
  INVX2 U1694 ( .A(n835), .Y(n1330) );
  MUX2X1 U1695 ( .B(core_block[246]), .A(n2148), .S(n2174), .Y(n836) );
  INVX2 U1696 ( .A(n836), .Y(n1329) );
  MUX2X1 U1697 ( .B(core_block[245]), .A(n2146), .S(n2174), .Y(n837) );
  INVX2 U1698 ( .A(n837), .Y(n1328) );
  MUX2X1 U1699 ( .B(core_block[244]), .A(n2144), .S(n2174), .Y(n838) );
  INVX2 U1700 ( .A(n838), .Y(n1327) );
  MUX2X1 U1701 ( .B(core_block[243]), .A(n2142), .S(n2174), .Y(n839) );
  INVX2 U1702 ( .A(n839), .Y(n1326) );
  MUX2X1 U1703 ( .B(core_block[242]), .A(n2140), .S(n2174), .Y(n840) );
  INVX2 U1704 ( .A(n840), .Y(n1325) );
  MUX2X1 U1705 ( .B(core_block[241]), .A(n2138), .S(n2174), .Y(n841) );
  INVX2 U1706 ( .A(n841), .Y(n1324) );
  MUX2X1 U1707 ( .B(core_block[240]), .A(n2136), .S(n2174), .Y(n842) );
  INVX2 U1708 ( .A(n842), .Y(n1323) );
  MUX2X1 U1709 ( .B(core_block[239]), .A(n2134), .S(n2174), .Y(n843) );
  INVX2 U1710 ( .A(n843), .Y(n1322) );
  MUX2X1 U1711 ( .B(core_block[238]), .A(n2132), .S(n2174), .Y(n844) );
  INVX2 U1712 ( .A(n844), .Y(n1321) );
  MUX2X1 U1713 ( .B(core_block[237]), .A(n2130), .S(n2174), .Y(n845) );
  INVX2 U1714 ( .A(n845), .Y(n1320) );
  MUX2X1 U1715 ( .B(core_block[236]), .A(n2128), .S(n2174), .Y(n846) );
  INVX2 U1716 ( .A(n846), .Y(n1319) );
  MUX2X1 U1717 ( .B(core_block[235]), .A(n2126), .S(n2174), .Y(n847) );
  INVX2 U1718 ( .A(n847), .Y(n1318) );
  MUX2X1 U1719 ( .B(core_block[234]), .A(n2124), .S(n2174), .Y(n848) );
  INVX2 U1720 ( .A(n848), .Y(n1317) );
  MUX2X1 U1721 ( .B(core_block[233]), .A(n2122), .S(n2174), .Y(n849) );
  INVX2 U1722 ( .A(n849), .Y(n1316) );
  MUX2X1 U1723 ( .B(core_block[232]), .A(n2120), .S(n2174), .Y(n850) );
  INVX2 U1724 ( .A(n850), .Y(n1315) );
  MUX2X1 U1725 ( .B(core_block[231]), .A(n2118), .S(n2174), .Y(n851) );
  INVX2 U1726 ( .A(n851), .Y(n1314) );
  MUX2X1 U1727 ( .B(core_block[230]), .A(n2116), .S(n2174), .Y(n852) );
  INVX2 U1728 ( .A(n852), .Y(n1313) );
  MUX2X1 U1729 ( .B(core_block[229]), .A(n2114), .S(n2174), .Y(n853) );
  INVX2 U1730 ( .A(n853), .Y(n1312) );
  MUX2X1 U1731 ( .B(core_block[228]), .A(n2112), .S(n2174), .Y(n854) );
  INVX2 U1732 ( .A(n854), .Y(n1311) );
  MUX2X1 U1733 ( .B(core_block[227]), .A(n2110), .S(n2174), .Y(n855) );
  INVX2 U1734 ( .A(n855), .Y(n1310) );
  MUX2X1 U1735 ( .B(core_block[226]), .A(n2108), .S(n2174), .Y(n856) );
  INVX2 U1736 ( .A(n856), .Y(n1309) );
  MUX2X1 U1737 ( .B(core_block[225]), .A(n2172), .S(n2174), .Y(n857) );
  INVX2 U1738 ( .A(n857), .Y(n1308) );
  MUX2X1 U1739 ( .B(core_block[224]), .A(n2170), .S(n2174), .Y(n858) );
  INVX2 U1740 ( .A(n858), .Y(n1307) );
  MUX2X1 U1741 ( .B(core_block[223]), .A(n2166), .S(n2236), .Y(n859) );
  INVX2 U1742 ( .A(n859), .Y(n1306) );
  MUX2X1 U1743 ( .B(core_block[222]), .A(n2164), .S(n2236), .Y(n860) );
  INVX2 U1744 ( .A(n860), .Y(n1305) );
  MUX2X1 U1745 ( .B(core_block[221]), .A(n2162), .S(n2236), .Y(n861) );
  INVX2 U1746 ( .A(n861), .Y(n1304) );
  MUX2X1 U1747 ( .B(core_block[220]), .A(n2160), .S(n2236), .Y(n862) );
  INVX2 U1748 ( .A(n862), .Y(n1303) );
  MUX2X1 U1749 ( .B(core_block[219]), .A(n2158), .S(n2236), .Y(n863) );
  INVX2 U1750 ( .A(n863), .Y(n1302) );
  MUX2X1 U1751 ( .B(core_block[218]), .A(n2156), .S(n2236), .Y(n864) );
  INVX2 U1752 ( .A(n864), .Y(n1301) );
  MUX2X1 U1753 ( .B(core_block[217]), .A(n2154), .S(n2236), .Y(n865) );
  INVX2 U1754 ( .A(n865), .Y(n1300) );
  MUX2X1 U1755 ( .B(core_block[216]), .A(n2152), .S(n2236), .Y(n866) );
  INVX2 U1756 ( .A(n866), .Y(n1299) );
  MUX2X1 U1757 ( .B(core_block[215]), .A(n2150), .S(n2236), .Y(n867) );
  INVX2 U1758 ( .A(n867), .Y(n1298) );
  MUX2X1 U1759 ( .B(core_block[214]), .A(n2148), .S(n2236), .Y(n868) );
  INVX2 U1760 ( .A(n868), .Y(n1297) );
  MUX2X1 U1761 ( .B(core_block[213]), .A(n2146), .S(n2236), .Y(n869) );
  INVX2 U1762 ( .A(n869), .Y(n1296) );
  MUX2X1 U1763 ( .B(core_block[212]), .A(n2144), .S(n2236), .Y(n870) );
  INVX2 U1764 ( .A(n870), .Y(n1295) );
  MUX2X1 U1765 ( .B(core_block[211]), .A(n2142), .S(n2236), .Y(n871) );
  INVX2 U1766 ( .A(n871), .Y(n1294) );
  MUX2X1 U1767 ( .B(core_block[210]), .A(n2140), .S(n2236), .Y(n872) );
  INVX2 U1768 ( .A(n872), .Y(n1293) );
  MUX2X1 U1769 ( .B(core_block[209]), .A(n2138), .S(n2236), .Y(n873) );
  INVX2 U1770 ( .A(n873), .Y(n1292) );
  MUX2X1 U1771 ( .B(core_block[208]), .A(n2136), .S(n2236), .Y(n874) );
  INVX2 U1772 ( .A(n874), .Y(n1291) );
  MUX2X1 U1773 ( .B(core_block[207]), .A(n2134), .S(n2236), .Y(n875) );
  INVX2 U1774 ( .A(n875), .Y(n1290) );
  MUX2X1 U1775 ( .B(core_block[206]), .A(n2132), .S(n2236), .Y(n876) );
  INVX2 U1776 ( .A(n876), .Y(n1289) );
  MUX2X1 U1777 ( .B(core_block[205]), .A(n2130), .S(n2236), .Y(n877) );
  INVX2 U1778 ( .A(n877), .Y(n1288) );
  MUX2X1 U1779 ( .B(core_block[204]), .A(n2128), .S(n2236), .Y(n878) );
  INVX2 U1780 ( .A(n878), .Y(n1287) );
  MUX2X1 U1781 ( .B(core_block[203]), .A(n2126), .S(n2236), .Y(n879) );
  INVX2 U1782 ( .A(n879), .Y(n1286) );
  MUX2X1 U1783 ( .B(core_block[202]), .A(n2124), .S(n2236), .Y(n880) );
  INVX2 U1784 ( .A(n880), .Y(n1285) );
  MUX2X1 U1785 ( .B(core_block[201]), .A(n2122), .S(n2236), .Y(n881) );
  INVX2 U1786 ( .A(n881), .Y(n1284) );
  MUX2X1 U1787 ( .B(core_block[200]), .A(n2120), .S(n2236), .Y(n882) );
  INVX2 U1788 ( .A(n882), .Y(n1283) );
  MUX2X1 U1789 ( .B(core_block[199]), .A(n2118), .S(n2236), .Y(n883) );
  INVX2 U1790 ( .A(n883), .Y(n1282) );
  MUX2X1 U1791 ( .B(core_block[198]), .A(n2116), .S(n2236), .Y(n884) );
  INVX2 U1792 ( .A(n884), .Y(n1281) );
  MUX2X1 U1793 ( .B(core_block[197]), .A(n2114), .S(n2236), .Y(n885) );
  INVX2 U1794 ( .A(n885), .Y(n1280) );
  MUX2X1 U1795 ( .B(core_block[196]), .A(n2112), .S(n2236), .Y(n886) );
  INVX2 U1796 ( .A(n886), .Y(n1279) );
  MUX2X1 U1797 ( .B(core_block[195]), .A(n2110), .S(n2236), .Y(n887) );
  INVX2 U1798 ( .A(n887), .Y(n1278) );
  MUX2X1 U1799 ( .B(core_block[194]), .A(n2108), .S(n2236), .Y(n888) );
  INVX2 U1800 ( .A(n888), .Y(n1277) );
  MUX2X1 U1801 ( .B(core_block[193]), .A(n2172), .S(n2236), .Y(n889) );
  INVX2 U1802 ( .A(n889), .Y(n1276) );
  MUX2X1 U1803 ( .B(core_block[192]), .A(n2170), .S(n2236), .Y(n890) );
  INVX2 U1804 ( .A(n890), .Y(n1275) );
  MUX2X1 U1805 ( .B(core_block[191]), .A(n2166), .S(n2234), .Y(n891) );
  INVX2 U1806 ( .A(n891), .Y(n1274) );
  MUX2X1 U1807 ( .B(core_block[190]), .A(n2164), .S(n2234), .Y(n892) );
  INVX2 U1808 ( .A(n892), .Y(n1273) );
  MUX2X1 U1809 ( .B(core_block[189]), .A(n2162), .S(n2234), .Y(n893) );
  INVX2 U1810 ( .A(n893), .Y(n1272) );
  MUX2X1 U1811 ( .B(core_block[188]), .A(n2160), .S(n2234), .Y(n894) );
  INVX2 U1812 ( .A(n894), .Y(n1271) );
  MUX2X1 U1813 ( .B(core_block[187]), .A(n2158), .S(n2234), .Y(n895) );
  INVX2 U1814 ( .A(n895), .Y(n1270) );
  MUX2X1 U1815 ( .B(core_block[186]), .A(n2156), .S(n2234), .Y(n896) );
  INVX2 U1816 ( .A(n896), .Y(n1269) );
  MUX2X1 U1817 ( .B(core_block[185]), .A(n2154), .S(n2234), .Y(n897) );
  INVX2 U1818 ( .A(n897), .Y(n1268) );
  MUX2X1 U1819 ( .B(core_block[184]), .A(n2152), .S(n2234), .Y(n898) );
  INVX2 U1820 ( .A(n898), .Y(n1267) );
  MUX2X1 U1821 ( .B(core_block[183]), .A(n2150), .S(n2234), .Y(n899) );
  INVX2 U1822 ( .A(n899), .Y(n1266) );
  MUX2X1 U1823 ( .B(core_block[182]), .A(n2148), .S(n2234), .Y(n900) );
  INVX2 U1824 ( .A(n900), .Y(n1265) );
  MUX2X1 U1825 ( .B(core_block[181]), .A(n2146), .S(n2234), .Y(n901) );
  INVX2 U1826 ( .A(n901), .Y(n1264) );
  MUX2X1 U1827 ( .B(core_block[180]), .A(n2144), .S(n2234), .Y(n902) );
  INVX2 U1828 ( .A(n902), .Y(n1263) );
  MUX2X1 U1829 ( .B(core_block[179]), .A(n2142), .S(n2234), .Y(n903) );
  INVX2 U1830 ( .A(n903), .Y(n1262) );
  MUX2X1 U1831 ( .B(core_block[178]), .A(n2140), .S(n2234), .Y(n904) );
  INVX2 U1832 ( .A(n904), .Y(n1261) );
  MUX2X1 U1833 ( .B(core_block[177]), .A(n2138), .S(n2234), .Y(n905) );
  INVX2 U1834 ( .A(n905), .Y(n1260) );
  MUX2X1 U1835 ( .B(core_block[176]), .A(n2136), .S(n2234), .Y(n906) );
  INVX2 U1836 ( .A(n906), .Y(n1259) );
  MUX2X1 U1837 ( .B(core_block[175]), .A(n2134), .S(n2234), .Y(n907) );
  INVX2 U1838 ( .A(n907), .Y(n1258) );
  MUX2X1 U1839 ( .B(core_block[174]), .A(n2132), .S(n2234), .Y(n908) );
  INVX2 U1840 ( .A(n908), .Y(n1257) );
  MUX2X1 U1841 ( .B(core_block[173]), .A(n2130), .S(n2234), .Y(n909) );
  INVX2 U1842 ( .A(n909), .Y(n1256) );
  MUX2X1 U1843 ( .B(core_block[172]), .A(n2128), .S(n2234), .Y(n910) );
  INVX2 U1844 ( .A(n910), .Y(n1255) );
  MUX2X1 U1845 ( .B(core_block[171]), .A(n2126), .S(n2234), .Y(n911) );
  INVX2 U1846 ( .A(n911), .Y(n1254) );
  MUX2X1 U1847 ( .B(core_block[170]), .A(n2124), .S(n2234), .Y(n912) );
  INVX2 U1848 ( .A(n912), .Y(n1253) );
  MUX2X1 U1849 ( .B(core_block[169]), .A(n2122), .S(n2234), .Y(n913) );
  INVX2 U1850 ( .A(n913), .Y(n1252) );
  MUX2X1 U1851 ( .B(core_block[168]), .A(n2120), .S(n2234), .Y(n914) );
  INVX2 U1852 ( .A(n914), .Y(n1251) );
  MUX2X1 U1853 ( .B(core_block[167]), .A(n2118), .S(n2234), .Y(n915) );
  INVX2 U1854 ( .A(n915), .Y(n1250) );
  MUX2X1 U1855 ( .B(core_block[166]), .A(n2116), .S(n2234), .Y(n916) );
  INVX2 U1856 ( .A(n916), .Y(n1249) );
  MUX2X1 U1857 ( .B(core_block[165]), .A(n2114), .S(n2234), .Y(n917) );
  INVX2 U1858 ( .A(n917), .Y(n1248) );
  MUX2X1 U1859 ( .B(core_block[164]), .A(n2112), .S(n2234), .Y(n918) );
  INVX2 U1860 ( .A(n918), .Y(n1247) );
  MUX2X1 U1861 ( .B(core_block[163]), .A(n2110), .S(n2234), .Y(n919) );
  INVX2 U1862 ( .A(n919), .Y(n1246) );
  MUX2X1 U1863 ( .B(core_block[162]), .A(n2108), .S(n2234), .Y(n920) );
  INVX2 U1864 ( .A(n920), .Y(n1245) );
  MUX2X1 U1865 ( .B(core_block[161]), .A(n2172), .S(n2234), .Y(n921) );
  INVX2 U1866 ( .A(n921), .Y(n1244) );
  MUX2X1 U1867 ( .B(core_block[160]), .A(n2170), .S(n2234), .Y(n922) );
  INVX2 U1868 ( .A(n922), .Y(n1243) );
  MUX2X1 U1869 ( .B(core_block[159]), .A(n2166), .S(n2232), .Y(n923) );
  INVX2 U1870 ( .A(n923), .Y(n1242) );
  MUX2X1 U1871 ( .B(core_block[158]), .A(n2164), .S(n2232), .Y(n924) );
  INVX2 U1872 ( .A(n924), .Y(n1241) );
  MUX2X1 U1873 ( .B(core_block[157]), .A(n2162), .S(n2232), .Y(n925) );
  INVX2 U1874 ( .A(n925), .Y(n1240) );
  MUX2X1 U1875 ( .B(core_block[156]), .A(n2160), .S(n2232), .Y(n926) );
  INVX2 U1876 ( .A(n926), .Y(n1239) );
  MUX2X1 U1877 ( .B(core_block[155]), .A(n2158), .S(n2232), .Y(n927) );
  INVX2 U1878 ( .A(n927), .Y(n1238) );
  MUX2X1 U1879 ( .B(core_block[154]), .A(n2156), .S(n2232), .Y(n928) );
  INVX2 U1880 ( .A(n928), .Y(n1237) );
  MUX2X1 U1881 ( .B(core_block[153]), .A(n2154), .S(n2232), .Y(n929) );
  INVX2 U1882 ( .A(n929), .Y(n1236) );
  MUX2X1 U1883 ( .B(core_block[152]), .A(n2152), .S(n2232), .Y(n930) );
  INVX2 U1884 ( .A(n930), .Y(n1235) );
  MUX2X1 U1885 ( .B(core_block[151]), .A(n2150), .S(n2232), .Y(n931) );
  INVX2 U1886 ( .A(n931), .Y(n1234) );
  MUX2X1 U1887 ( .B(core_block[150]), .A(n2148), .S(n2232), .Y(n932) );
  INVX2 U1888 ( .A(n932), .Y(n1233) );
  MUX2X1 U1889 ( .B(core_block[149]), .A(n2146), .S(n2232), .Y(n933) );
  INVX2 U1890 ( .A(n933), .Y(n1232) );
  MUX2X1 U1891 ( .B(core_block[148]), .A(n2144), .S(n2232), .Y(n934) );
  INVX2 U1892 ( .A(n934), .Y(n1231) );
  MUX2X1 U1893 ( .B(core_block[147]), .A(n2142), .S(n2232), .Y(n935) );
  INVX2 U1894 ( .A(n935), .Y(n1230) );
  MUX2X1 U1895 ( .B(core_block[146]), .A(n2140), .S(n2232), .Y(n936) );
  INVX2 U1896 ( .A(n936), .Y(n1229) );
  MUX2X1 U1897 ( .B(core_block[145]), .A(n2138), .S(n2232), .Y(n937) );
  INVX2 U1898 ( .A(n937), .Y(n1228) );
  MUX2X1 U1899 ( .B(core_block[144]), .A(n2136), .S(n2232), .Y(n938) );
  INVX2 U1900 ( .A(n938), .Y(n1227) );
  MUX2X1 U1901 ( .B(core_block[143]), .A(n2134), .S(n2232), .Y(n939) );
  INVX2 U1902 ( .A(n939), .Y(n1226) );
  MUX2X1 U1903 ( .B(core_block[142]), .A(n2132), .S(n2232), .Y(n940) );
  INVX2 U1904 ( .A(n940), .Y(n1225) );
  MUX2X1 U1905 ( .B(core_block[141]), .A(n2130), .S(n2232), .Y(n941) );
  INVX2 U1906 ( .A(n941), .Y(n1224) );
  MUX2X1 U1907 ( .B(core_block[140]), .A(n2128), .S(n2232), .Y(n942) );
  INVX2 U1908 ( .A(n942), .Y(n1223) );
  MUX2X1 U1909 ( .B(core_block[139]), .A(n2126), .S(n2232), .Y(n943) );
  INVX2 U1910 ( .A(n943), .Y(n1222) );
  MUX2X1 U1911 ( .B(core_block[138]), .A(n2124), .S(n2232), .Y(n944) );
  INVX2 U1912 ( .A(n944), .Y(n1221) );
  MUX2X1 U1913 ( .B(core_block[137]), .A(n2122), .S(n2232), .Y(n945) );
  INVX2 U1914 ( .A(n945), .Y(n1220) );
  MUX2X1 U1915 ( .B(core_block[136]), .A(n2120), .S(n2232), .Y(n946) );
  INVX2 U1916 ( .A(n946), .Y(n1219) );
  MUX2X1 U1917 ( .B(core_block[135]), .A(n2118), .S(n2232), .Y(n947) );
  INVX2 U1918 ( .A(n947), .Y(n1218) );
  MUX2X1 U1919 ( .B(core_block[134]), .A(n2116), .S(n2232), .Y(n948) );
  INVX2 U1920 ( .A(n948), .Y(n1217) );
  MUX2X1 U1921 ( .B(core_block[133]), .A(n2114), .S(n2232), .Y(n949) );
  INVX2 U1922 ( .A(n949), .Y(n1216) );
  MUX2X1 U1923 ( .B(core_block[132]), .A(n2112), .S(n2232), .Y(n950) );
  INVX2 U1924 ( .A(n950), .Y(n1215) );
  MUX2X1 U1925 ( .B(core_block[131]), .A(n2110), .S(n2232), .Y(n951) );
  INVX2 U1926 ( .A(n951), .Y(n1214) );
  MUX2X1 U1927 ( .B(core_block[130]), .A(n2108), .S(n2232), .Y(n952) );
  INVX2 U1928 ( .A(n952), .Y(n1213) );
  MUX2X1 U1929 ( .B(core_block[129]), .A(n2172), .S(n2232), .Y(n953) );
  INVX2 U1930 ( .A(n953), .Y(n1212) );
  MUX2X1 U1931 ( .B(core_block[128]), .A(n2170), .S(n2232), .Y(n954) );
  INVX2 U1932 ( .A(n954), .Y(n1211) );
  MUX2X1 U1933 ( .B(core_block[127]), .A(n2166), .S(n2230), .Y(n955) );
  INVX2 U1934 ( .A(n955), .Y(n1210) );
  MUX2X1 U1935 ( .B(core_block[126]), .A(n2164), .S(n2230), .Y(n956) );
  INVX2 U1936 ( .A(n956), .Y(n1209) );
  MUX2X1 U1937 ( .B(core_block[125]), .A(n2162), .S(n2230), .Y(n957) );
  INVX2 U1938 ( .A(n957), .Y(n1208) );
  MUX2X1 U1939 ( .B(core_block[124]), .A(n2160), .S(n2230), .Y(n958) );
  INVX2 U1940 ( .A(n958), .Y(n1207) );
  MUX2X1 U1941 ( .B(core_block[123]), .A(n2158), .S(n2230), .Y(n959) );
  INVX2 U1942 ( .A(n959), .Y(n1206) );
  MUX2X1 U1943 ( .B(core_block[122]), .A(n2156), .S(n2230), .Y(n960) );
  INVX2 U1944 ( .A(n960), .Y(n1205) );
  MUX2X1 U1945 ( .B(core_block[121]), .A(n2154), .S(n2230), .Y(n961) );
  INVX2 U1946 ( .A(n961), .Y(n1204) );
  MUX2X1 U1947 ( .B(core_block[120]), .A(n2152), .S(n2230), .Y(n962) );
  INVX2 U1948 ( .A(n962), .Y(n1203) );
  MUX2X1 U1949 ( .B(core_block[119]), .A(n2150), .S(n2230), .Y(n963) );
  INVX2 U1950 ( .A(n963), .Y(n1202) );
  MUX2X1 U1951 ( .B(core_block[118]), .A(n2148), .S(n2230), .Y(n964) );
  INVX2 U1952 ( .A(n964), .Y(n1201) );
  MUX2X1 U1953 ( .B(core_block[117]), .A(n2146), .S(n2230), .Y(n965) );
  INVX2 U1954 ( .A(n965), .Y(n1200) );
  MUX2X1 U1955 ( .B(core_block[116]), .A(n2144), .S(n2230), .Y(n966) );
  INVX2 U1956 ( .A(n966), .Y(n1199) );
  MUX2X1 U1957 ( .B(core_block[115]), .A(n2142), .S(n2230), .Y(n967) );
  INVX2 U1958 ( .A(n967), .Y(n1198) );
  MUX2X1 U1959 ( .B(core_block[114]), .A(n2140), .S(n2230), .Y(n968) );
  INVX2 U1960 ( .A(n968), .Y(n1197) );
  MUX2X1 U1961 ( .B(core_block[113]), .A(n2138), .S(n2230), .Y(n969) );
  INVX2 U1962 ( .A(n969), .Y(n1196) );
  MUX2X1 U1963 ( .B(core_block[112]), .A(n2136), .S(n2230), .Y(n970) );
  INVX2 U1964 ( .A(n970), .Y(n1195) );
  MUX2X1 U1965 ( .B(core_block[111]), .A(n2134), .S(n2230), .Y(n971) );
  INVX2 U1966 ( .A(n971), .Y(n1194) );
  MUX2X1 U1967 ( .B(core_block[110]), .A(n2132), .S(n2230), .Y(n972) );
  INVX2 U1968 ( .A(n972), .Y(n1193) );
  MUX2X1 U1969 ( .B(core_block[109]), .A(n2130), .S(n2230), .Y(n973) );
  INVX2 U1970 ( .A(n973), .Y(n1192) );
  MUX2X1 U1971 ( .B(core_block[108]), .A(n2128), .S(n2230), .Y(n974) );
  INVX2 U1972 ( .A(n974), .Y(n1191) );
  MUX2X1 U1973 ( .B(core_block[107]), .A(n2126), .S(n2230), .Y(n975) );
  INVX2 U1974 ( .A(n975), .Y(n1190) );
  MUX2X1 U1975 ( .B(core_block[106]), .A(n2124), .S(n2230), .Y(n976) );
  INVX2 U1976 ( .A(n976), .Y(n1189) );
  MUX2X1 U1977 ( .B(core_block[105]), .A(n2122), .S(n2230), .Y(n977) );
  INVX2 U1978 ( .A(n977), .Y(n1188) );
  MUX2X1 U1979 ( .B(core_block[104]), .A(n2120), .S(n2230), .Y(n978) );
  INVX2 U1980 ( .A(n978), .Y(n1187) );
  MUX2X1 U1981 ( .B(core_block[103]), .A(n2118), .S(n2230), .Y(n979) );
  INVX2 U1982 ( .A(n979), .Y(n1186) );
  MUX2X1 U1983 ( .B(core_block[102]), .A(n2116), .S(n2230), .Y(n980) );
  INVX2 U1984 ( .A(n980), .Y(n1185) );
  MUX2X1 U1985 ( .B(core_block[101]), .A(n2114), .S(n2230), .Y(n981) );
  INVX2 U1986 ( .A(n981), .Y(n1184) );
  MUX2X1 U1987 ( .B(core_block[100]), .A(n2112), .S(n2230), .Y(n982) );
  INVX2 U1988 ( .A(n982), .Y(n1183) );
  MUX2X1 U1989 ( .B(core_block[99]), .A(n2110), .S(n2230), .Y(n983) );
  INVX2 U1990 ( .A(n983), .Y(n1182) );
  MUX2X1 U1991 ( .B(core_block[98]), .A(n2108), .S(n2230), .Y(n984) );
  INVX2 U1992 ( .A(n984), .Y(n1181) );
  MUX2X1 U1993 ( .B(core_block[97]), .A(n2172), .S(n2230), .Y(n985) );
  INVX2 U1994 ( .A(n985), .Y(n1180) );
  MUX2X1 U1995 ( .B(core_block[96]), .A(n2170), .S(n2230), .Y(n986) );
  INVX2 U1996 ( .A(n986), .Y(n1179) );
  MUX2X1 U1997 ( .B(core_block[95]), .A(n2166), .S(n2228), .Y(n987) );
  INVX2 U1998 ( .A(n987), .Y(n1178) );
  MUX2X1 U1999 ( .B(core_block[94]), .A(n2164), .S(n2228), .Y(n988) );
  INVX2 U2000 ( .A(n988), .Y(n1177) );
  MUX2X1 U2001 ( .B(core_block[93]), .A(n2162), .S(n2228), .Y(n989) );
  INVX2 U2002 ( .A(n989), .Y(n1176) );
  MUX2X1 U2003 ( .B(core_block[92]), .A(n2160), .S(n2228), .Y(n990) );
  INVX2 U2004 ( .A(n990), .Y(n1175) );
  MUX2X1 U2005 ( .B(core_block[91]), .A(n2158), .S(n2228), .Y(n991) );
  INVX2 U2006 ( .A(n991), .Y(n1174) );
  MUX2X1 U2007 ( .B(core_block[90]), .A(n2156), .S(n2228), .Y(n992) );
  INVX2 U2008 ( .A(n992), .Y(n1173) );
  MUX2X1 U2009 ( .B(core_block[89]), .A(n2154), .S(n2228), .Y(n993) );
  INVX2 U2010 ( .A(n993), .Y(n1172) );
  MUX2X1 U2011 ( .B(core_block[88]), .A(n2152), .S(n2228), .Y(n994) );
  INVX2 U2012 ( .A(n994), .Y(n1171) );
  MUX2X1 U2013 ( .B(core_block[87]), .A(n2150), .S(n2228), .Y(n995) );
  INVX2 U2014 ( .A(n995), .Y(n1170) );
  MUX2X1 U2015 ( .B(core_block[86]), .A(n2148), .S(n2228), .Y(n996) );
  INVX2 U2016 ( .A(n996), .Y(n1169) );
  MUX2X1 U2017 ( .B(core_block[85]), .A(n2146), .S(n2228), .Y(n997) );
  INVX2 U2018 ( .A(n997), .Y(n1168) );
  MUX2X1 U2019 ( .B(core_block[84]), .A(n2144), .S(n2228), .Y(n998) );
  INVX2 U2020 ( .A(n998), .Y(n1167) );
  MUX2X1 U2021 ( .B(core_block[83]), .A(n2142), .S(n2228), .Y(n999) );
  INVX2 U2022 ( .A(n999), .Y(n1166) );
  MUX2X1 U2023 ( .B(core_block[82]), .A(n2140), .S(n2228), .Y(n1000) );
  INVX2 U2024 ( .A(n1000), .Y(n1165) );
  MUX2X1 U2025 ( .B(core_block[81]), .A(n2138), .S(n2228), .Y(n1001) );
  INVX2 U2026 ( .A(n1001), .Y(n1164) );
  MUX2X1 U2027 ( .B(core_block[80]), .A(n2136), .S(n2228), .Y(n1002) );
  INVX2 U2028 ( .A(n1002), .Y(n1163) );
  MUX2X1 U2029 ( .B(core_block[79]), .A(n2134), .S(n2228), .Y(n1003) );
  INVX2 U2030 ( .A(n1003), .Y(n1162) );
  MUX2X1 U2031 ( .B(core_block[78]), .A(n2132), .S(n2228), .Y(n1004) );
  INVX2 U2032 ( .A(n1004), .Y(n1161) );
  MUX2X1 U2033 ( .B(core_block[77]), .A(n2130), .S(n2228), .Y(n1005) );
  INVX2 U2034 ( .A(n1005), .Y(n1160) );
  MUX2X1 U2035 ( .B(core_block[76]), .A(n2128), .S(n2228), .Y(n1006) );
  INVX2 U2036 ( .A(n1006), .Y(n1159) );
  MUX2X1 U2037 ( .B(core_block[75]), .A(n2126), .S(n2228), .Y(n1007) );
  INVX2 U2038 ( .A(n1007), .Y(n1158) );
  MUX2X1 U2039 ( .B(core_block[74]), .A(n2124), .S(n2228), .Y(n1008) );
  INVX2 U2040 ( .A(n1008), .Y(n1157) );
  MUX2X1 U2041 ( .B(core_block[73]), .A(n2122), .S(n2228), .Y(n1009) );
  INVX2 U2042 ( .A(n1009), .Y(n1156) );
  MUX2X1 U2043 ( .B(core_block[72]), .A(n2120), .S(n2228), .Y(n1010) );
  INVX2 U2044 ( .A(n1010), .Y(n1155) );
  MUX2X1 U2045 ( .B(core_block[71]), .A(n2118), .S(n2228), .Y(n1011) );
  INVX2 U2046 ( .A(n1011), .Y(n1154) );
  MUX2X1 U2047 ( .B(core_block[70]), .A(n2116), .S(n2228), .Y(n1012) );
  INVX2 U2048 ( .A(n1012), .Y(n1153) );
  MUX2X1 U2049 ( .B(core_block[69]), .A(n2114), .S(n2228), .Y(n1013) );
  INVX2 U2050 ( .A(n1013), .Y(n1152) );
  MUX2X1 U2051 ( .B(core_block[68]), .A(n2112), .S(n2228), .Y(n1014) );
  INVX2 U2052 ( .A(n1014), .Y(n1151) );
  MUX2X1 U2053 ( .B(core_block[67]), .A(n2110), .S(n2228), .Y(n1015) );
  INVX2 U2054 ( .A(n1015), .Y(n1150) );
  MUX2X1 U2055 ( .B(core_block[66]), .A(n2108), .S(n2228), .Y(n1016) );
  INVX2 U2056 ( .A(n1016), .Y(n1149) );
  MUX2X1 U2057 ( .B(core_block[65]), .A(n2172), .S(n2228), .Y(n1017) );
  INVX2 U2058 ( .A(n1017), .Y(n1148) );
  MUX2X1 U2059 ( .B(core_block[64]), .A(n2170), .S(n2228), .Y(n1018) );
  INVX2 U2060 ( .A(n1018), .Y(n1147) );
  MUX2X1 U2061 ( .B(core_block[63]), .A(n2166), .S(n2226), .Y(n1019) );
  INVX2 U2062 ( .A(n1019), .Y(n1146) );
  MUX2X1 U2063 ( .B(core_block[62]), .A(n2164), .S(n2226), .Y(n1020) );
  INVX2 U2064 ( .A(n1020), .Y(n1145) );
  MUX2X1 U2065 ( .B(core_block[61]), .A(n2162), .S(n2226), .Y(n1021) );
  INVX2 U2066 ( .A(n1021), .Y(n1144) );
  MUX2X1 U2067 ( .B(core_block[60]), .A(n2160), .S(n2226), .Y(n1022) );
  INVX2 U2068 ( .A(n1022), .Y(n1143) );
  MUX2X1 U2069 ( .B(core_block[59]), .A(n2158), .S(n2226), .Y(n1023) );
  INVX2 U2070 ( .A(n1023), .Y(n1142) );
  MUX2X1 U2071 ( .B(core_block[58]), .A(n2156), .S(n2226), .Y(n1024) );
  INVX2 U2072 ( .A(n1024), .Y(n1141) );
  MUX2X1 U2073 ( .B(core_block[57]), .A(n2154), .S(n2226), .Y(n1025) );
  INVX2 U2074 ( .A(n1025), .Y(n1140) );
  MUX2X1 U2075 ( .B(core_block[56]), .A(n2152), .S(n2226), .Y(n1026) );
  INVX2 U2076 ( .A(n1026), .Y(n1139) );
  MUX2X1 U2077 ( .B(core_block[55]), .A(n2150), .S(n2226), .Y(n1027) );
  INVX2 U2078 ( .A(n1027), .Y(n1138) );
  MUX2X1 U2079 ( .B(core_block[54]), .A(n2148), .S(n2226), .Y(n1028) );
  INVX2 U2080 ( .A(n1028), .Y(n1137) );
  MUX2X1 U2081 ( .B(core_block[53]), .A(n2146), .S(n2226), .Y(n1029) );
  INVX2 U2082 ( .A(n1029), .Y(n1136) );
  MUX2X1 U2083 ( .B(core_block[52]), .A(n2144), .S(n2226), .Y(n1030) );
  INVX2 U2084 ( .A(n1030), .Y(n1135) );
  MUX2X1 U2085 ( .B(core_block[51]), .A(n2142), .S(n2226), .Y(n1031) );
  INVX2 U2086 ( .A(n1031), .Y(n1134) );
  MUX2X1 U2087 ( .B(core_block[50]), .A(n2140), .S(n2226), .Y(n1032) );
  INVX2 U2088 ( .A(n1032), .Y(n1133) );
  MUX2X1 U2089 ( .B(core_block[49]), .A(n2138), .S(n2226), .Y(n1033) );
  INVX2 U2090 ( .A(n1033), .Y(n1132) );
  MUX2X1 U2091 ( .B(core_block[48]), .A(n2136), .S(n2226), .Y(n1034) );
  INVX2 U2092 ( .A(n1034), .Y(n1131) );
  MUX2X1 U2093 ( .B(core_block[47]), .A(n2134), .S(n2226), .Y(n1035) );
  INVX2 U2094 ( .A(n1035), .Y(n1130) );
  MUX2X1 U2095 ( .B(core_block[46]), .A(n2132), .S(n2226), .Y(n1036) );
  INVX2 U2096 ( .A(n1036), .Y(n1129) );
  MUX2X1 U2097 ( .B(core_block[45]), .A(n2130), .S(n2226), .Y(n1037) );
  INVX2 U2098 ( .A(n1037), .Y(n1128) );
  MUX2X1 U2099 ( .B(core_block[44]), .A(n2128), .S(n2226), .Y(n1038) );
  INVX2 U2100 ( .A(n1038), .Y(n1127) );
  MUX2X1 U2101 ( .B(core_block[43]), .A(n2126), .S(n2226), .Y(n1039) );
  INVX2 U2102 ( .A(n1039), .Y(n1126) );
  MUX2X1 U2103 ( .B(core_block[42]), .A(n2124), .S(n2226), .Y(n1040) );
  INVX2 U2104 ( .A(n1040), .Y(n1125) );
  MUX2X1 U2105 ( .B(core_block[41]), .A(n2122), .S(n2226), .Y(n1041) );
  INVX2 U2106 ( .A(n1041), .Y(n1124) );
  MUX2X1 U2107 ( .B(core_block[40]), .A(n2120), .S(n2226), .Y(n1042) );
  INVX2 U2108 ( .A(n1042), .Y(n1123) );
  MUX2X1 U2109 ( .B(core_block[39]), .A(n2118), .S(n2226), .Y(n1043) );
  INVX2 U2110 ( .A(n1043), .Y(n1122) );
  MUX2X1 U2111 ( .B(core_block[38]), .A(n2116), .S(n2226), .Y(n1044) );
  INVX2 U2112 ( .A(n1044), .Y(n1121) );
  MUX2X1 U2113 ( .B(core_block[37]), .A(n2114), .S(n2226), .Y(n1045) );
  INVX2 U2114 ( .A(n1045), .Y(n1120) );
  MUX2X1 U2115 ( .B(core_block[36]), .A(n2112), .S(n2226), .Y(n1046) );
  INVX2 U2116 ( .A(n1046), .Y(n1119) );
  MUX2X1 U2117 ( .B(core_block[35]), .A(n2110), .S(n2226), .Y(n1047) );
  INVX2 U2118 ( .A(n1047), .Y(n1118) );
  MUX2X1 U2119 ( .B(core_block[34]), .A(n2108), .S(n2226), .Y(n1048) );
  INVX2 U2120 ( .A(n1048), .Y(n1117) );
  MUX2X1 U2121 ( .B(core_block[33]), .A(n2172), .S(n2226), .Y(n1049) );
  INVX2 U2122 ( .A(n1049), .Y(n1116) );
  MUX2X1 U2123 ( .B(core_block[32]), .A(n2170), .S(n2226), .Y(n1050) );
  INVX2 U2124 ( .A(n1050), .Y(n1115) );
  MUX2X1 U2125 ( .B(core_block[31]), .A(n2166), .S(n2224), .Y(n1051) );
  INVX2 U2126 ( .A(n1051), .Y(n1114) );
  MUX2X1 U2127 ( .B(core_block[30]), .A(n2164), .S(n2224), .Y(n1052) );
  INVX2 U2128 ( .A(n1052), .Y(n1113) );
  MUX2X1 U2129 ( .B(core_block[29]), .A(n2162), .S(n2224), .Y(n1053) );
  INVX2 U2130 ( .A(n1053), .Y(n1112) );
  MUX2X1 U2131 ( .B(core_block[28]), .A(n2160), .S(n2224), .Y(n1054) );
  INVX2 U2132 ( .A(n1054), .Y(n1111) );
  MUX2X1 U2133 ( .B(core_block[27]), .A(n2158), .S(n2224), .Y(n1055) );
  INVX2 U2134 ( .A(n1055), .Y(n1110) );
  MUX2X1 U2135 ( .B(core_block[26]), .A(n2156), .S(n2224), .Y(n1056) );
  INVX2 U2136 ( .A(n1056), .Y(n1109) );
  MUX2X1 U2137 ( .B(core_block[25]), .A(n2154), .S(n2224), .Y(n1057) );
  INVX2 U2138 ( .A(n1057), .Y(n1108) );
  MUX2X1 U2139 ( .B(core_block[24]), .A(n2152), .S(n2224), .Y(n1058) );
  INVX2 U2140 ( .A(n1058), .Y(n1107) );
  MUX2X1 U2141 ( .B(core_block[23]), .A(n2150), .S(n2224), .Y(n1059) );
  INVX2 U2142 ( .A(n1059), .Y(n1106) );
  MUX2X1 U2143 ( .B(core_block[22]), .A(n2148), .S(n2224), .Y(n1060) );
  INVX2 U2144 ( .A(n1060), .Y(n1105) );
  MUX2X1 U2145 ( .B(core_block[21]), .A(n2146), .S(n2224), .Y(n1061) );
  INVX2 U2146 ( .A(n1061), .Y(n1104) );
  MUX2X1 U2147 ( .B(core_block[20]), .A(n2144), .S(n2224), .Y(n1062) );
  INVX2 U2148 ( .A(n1062), .Y(n1103) );
  MUX2X1 U2149 ( .B(core_block[19]), .A(n2142), .S(n2224), .Y(n1063) );
  INVX2 U2150 ( .A(n1063), .Y(n1102) );
  MUX2X1 U2151 ( .B(core_block[18]), .A(n2140), .S(n2224), .Y(n1064) );
  INVX2 U2152 ( .A(n1064), .Y(n1101) );
  MUX2X1 U2153 ( .B(core_block[17]), .A(n2138), .S(n2224), .Y(n1065) );
  INVX2 U2154 ( .A(n1065), .Y(n1100) );
  MUX2X1 U2155 ( .B(core_block[16]), .A(n2136), .S(n2224), .Y(n1066) );
  INVX2 U2156 ( .A(n1066), .Y(n1099) );
  MUX2X1 U2157 ( .B(core_block[15]), .A(n2134), .S(n2224), .Y(n1067) );
  INVX2 U2158 ( .A(n1067), .Y(n1098) );
  MUX2X1 U2159 ( .B(core_block[14]), .A(n2132), .S(n2224), .Y(n1068) );
  INVX2 U2160 ( .A(n1068), .Y(n1097) );
  MUX2X1 U2161 ( .B(core_block[13]), .A(n2130), .S(n2224), .Y(n1069) );
  INVX2 U2162 ( .A(n1069), .Y(n1096) );
  MUX2X1 U2163 ( .B(core_block[12]), .A(n2128), .S(n2224), .Y(n1070) );
  INVX2 U2164 ( .A(n1070), .Y(n1095) );
  MUX2X1 U2165 ( .B(core_block[11]), .A(n2126), .S(n2224), .Y(n1071) );
  INVX2 U2166 ( .A(n1071), .Y(n1094) );
  MUX2X1 U2167 ( .B(core_block[10]), .A(n2124), .S(n2224), .Y(n1072) );
  INVX2 U2168 ( .A(n1072), .Y(n1093) );
  MUX2X1 U2169 ( .B(core_block[9]), .A(n2122), .S(n2224), .Y(n1073) );
  INVX2 U2170 ( .A(n1073), .Y(n1092) );
  MUX2X1 U2171 ( .B(core_block[8]), .A(n2120), .S(n2224), .Y(n1074) );
  INVX2 U2172 ( .A(n1074), .Y(n1091) );
  MUX2X1 U2173 ( .B(core_block[7]), .A(n2118), .S(n2224), .Y(n1075) );
  INVX2 U2174 ( .A(n1075), .Y(n1090) );
  MUX2X1 U2175 ( .B(core_block[6]), .A(n2116), .S(n2224), .Y(n1076) );
  INVX2 U2176 ( .A(n1076), .Y(n1089) );
  MUX2X1 U2177 ( .B(core_block[5]), .A(n2114), .S(n2224), .Y(n1077) );
  INVX2 U2178 ( .A(n1077), .Y(n1088) );
  MUX2X1 U2179 ( .B(core_block[4]), .A(n2112), .S(n2224), .Y(n1078) );
  INVX2 U2180 ( .A(n1078), .Y(n1087) );
  MUX2X1 U2181 ( .B(core_block[3]), .A(n2110), .S(n2224), .Y(n1079) );
  INVX2 U2182 ( .A(n1079), .Y(n1086) );
  MUX2X1 U2183 ( .B(core_block[2]), .A(n2108), .S(n2224), .Y(n1080) );
  INVX2 U2184 ( .A(n1080), .Y(n1085) );
  MUX2X1 U2185 ( .B(core_block[1]), .A(n2172), .S(n2224), .Y(n1081) );
  INVX2 U2186 ( .A(n1081), .Y(n1084) );
  MUX2X1 U2187 ( .B(core_block[0]), .A(n2170), .S(n2224), .Y(n1082) );
  INVX2 U2188 ( .A(n1082), .Y(n1083) );
  blake2_core core ( .clk(clk), .reset_n(reset_n), .init(core_init), .next(
        core_next), .final_block(1'b0), .block(core_block), .data_length({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ready(core_ready), 
        .digest_valid(core_digest_valid) );
  INVX1 U2189 ( .A(N64), .Y(n2107) );
  INVX4 U2190 ( .A(n2107), .Y(n2108) );
  INVX1 U2191 ( .A(N65), .Y(n2109) );
  INVX4 U2192 ( .A(n2109), .Y(n2110) );
  INVX1 U2193 ( .A(N66), .Y(n2111) );
  INVX4 U2194 ( .A(n2111), .Y(n2112) );
  INVX1 U2195 ( .A(N67), .Y(n2113) );
  INVX4 U2196 ( .A(n2113), .Y(n2114) );
  INVX1 U2197 ( .A(N68), .Y(n2115) );
  INVX4 U2198 ( .A(n2115), .Y(n2116) );
  INVX1 U2199 ( .A(N69), .Y(n2117) );
  INVX4 U2200 ( .A(n2117), .Y(n2118) );
  INVX1 U2201 ( .A(N70), .Y(n2119) );
  INVX4 U2202 ( .A(n2119), .Y(n2120) );
  INVX1 U2203 ( .A(N71), .Y(n2121) );
  INVX4 U2204 ( .A(n2121), .Y(n2122) );
  INVX1 U2205 ( .A(N72), .Y(n2123) );
  INVX4 U2206 ( .A(n2123), .Y(n2124) );
  INVX1 U2207 ( .A(N73), .Y(n2125) );
  INVX4 U2208 ( .A(n2125), .Y(n2126) );
  INVX1 U2209 ( .A(N74), .Y(n2127) );
  INVX4 U2210 ( .A(n2127), .Y(n2128) );
  INVX1 U2211 ( .A(N75), .Y(n2129) );
  INVX4 U2212 ( .A(n2129), .Y(n2130) );
  INVX1 U2213 ( .A(N76), .Y(n2131) );
  INVX4 U2214 ( .A(n2131), .Y(n2132) );
  INVX1 U2215 ( .A(N77), .Y(n2133) );
  INVX4 U2216 ( .A(n2133), .Y(n2134) );
  INVX1 U2217 ( .A(N78), .Y(n2135) );
  INVX4 U2218 ( .A(n2135), .Y(n2136) );
  INVX1 U2219 ( .A(N79), .Y(n2137) );
  INVX4 U2220 ( .A(n2137), .Y(n2138) );
  INVX1 U2221 ( .A(N80), .Y(n2139) );
  INVX4 U2222 ( .A(n2139), .Y(n2140) );
  INVX1 U2223 ( .A(N81), .Y(n2141) );
  INVX4 U2224 ( .A(n2141), .Y(n2142) );
  INVX1 U2225 ( .A(N82), .Y(n2143) );
  INVX4 U2226 ( .A(n2143), .Y(n2144) );
  INVX1 U2227 ( .A(N83), .Y(n2145) );
  INVX4 U2228 ( .A(n2145), .Y(n2146) );
  INVX1 U2229 ( .A(N84), .Y(n2147) );
  INVX4 U2230 ( .A(n2147), .Y(n2148) );
  INVX1 U2231 ( .A(N85), .Y(n2149) );
  INVX4 U2232 ( .A(n2149), .Y(n2150) );
  INVX1 U2233 ( .A(N86), .Y(n2151) );
  INVX4 U2234 ( .A(n2151), .Y(n2152) );
  INVX1 U2235 ( .A(N87), .Y(n2153) );
  INVX4 U2236 ( .A(n2153), .Y(n2154) );
  INVX1 U2237 ( .A(N88), .Y(n2155) );
  INVX4 U2238 ( .A(n2155), .Y(n2156) );
  INVX1 U2239 ( .A(N89), .Y(n2157) );
  INVX4 U2240 ( .A(n2157), .Y(n2158) );
  INVX1 U2241 ( .A(N90), .Y(n2159) );
  INVX4 U2242 ( .A(n2159), .Y(n2160) );
  INVX1 U2243 ( .A(N91), .Y(n2161) );
  INVX4 U2244 ( .A(n2161), .Y(n2162) );
  INVX1 U2245 ( .A(N92), .Y(n2163) );
  INVX4 U2246 ( .A(n2163), .Y(n2164) );
  INVX1 U2247 ( .A(N93), .Y(n2165) );
  INVX4 U2248 ( .A(n2165), .Y(n2166) );
  INVX1 U2249 ( .A(n24), .Y(n2167) );
  INVX4 U2250 ( .A(n2167), .Y(n2168) );
  INVX1 U2251 ( .A(N59), .Y(n2169) );
  INVX4 U2252 ( .A(n2169), .Y(n2170) );
  INVX1 U2253 ( .A(N60), .Y(n2171) );
  INVX4 U2254 ( .A(n2171), .Y(n2172) );
  INVX1 U2255 ( .A(N100), .Y(n2173) );
  INVX4 U2256 ( .A(n2173), .Y(n2174) );
  INVX1 U2257 ( .A(N101), .Y(n2175) );
  INVX4 U2258 ( .A(n2175), .Y(n2176) );
  INVX1 U2259 ( .A(N102), .Y(n2177) );
  INVX4 U2260 ( .A(n2177), .Y(n2178) );
  INVX1 U2261 ( .A(N103), .Y(n2179) );
  INVX4 U2262 ( .A(n2179), .Y(n2180) );
  INVX1 U2263 ( .A(N104), .Y(n2181) );
  INVX4 U2264 ( .A(n2181), .Y(n2182) );
  INVX1 U2265 ( .A(N105), .Y(n2183) );
  INVX4 U2266 ( .A(n2183), .Y(n2184) );
  INVX1 U2267 ( .A(N106), .Y(n2185) );
  INVX4 U2268 ( .A(n2185), .Y(n2186) );
  INVX1 U2269 ( .A(N107), .Y(n2187) );
  INVX4 U2270 ( .A(n2187), .Y(n2188) );
  INVX1 U2271 ( .A(N108), .Y(n2189) );
  INVX4 U2272 ( .A(n2189), .Y(n2190) );
  INVX1 U2273 ( .A(N109), .Y(n2191) );
  INVX4 U2274 ( .A(n2191), .Y(n2192) );
  INVX1 U2275 ( .A(N110), .Y(n2193) );
  INVX4 U2276 ( .A(n2193), .Y(n2194) );
  INVX1 U2277 ( .A(N111), .Y(n2195) );
  INVX4 U2278 ( .A(n2195), .Y(n2196) );
  INVX1 U2279 ( .A(N112), .Y(n2197) );
  INVX4 U2280 ( .A(n2197), .Y(n2198) );
  INVX1 U2281 ( .A(N113), .Y(n2199) );
  INVX4 U2282 ( .A(n2199), .Y(n2200) );
  INVX1 U2283 ( .A(N114), .Y(n2201) );
  INVX4 U2284 ( .A(n2201), .Y(n2202) );
  INVX1 U2285 ( .A(N115), .Y(n2203) );
  INVX4 U2286 ( .A(n2203), .Y(n2204) );
  INVX1 U2287 ( .A(N116), .Y(n2205) );
  INVX4 U2288 ( .A(n2205), .Y(n2206) );
  INVX1 U2289 ( .A(N117), .Y(n2207) );
  INVX4 U2290 ( .A(n2207), .Y(n2208) );
  INVX1 U2291 ( .A(N118), .Y(n2209) );
  INVX4 U2292 ( .A(n2209), .Y(n2210) );
  INVX1 U2293 ( .A(N119), .Y(n2211) );
  INVX4 U2294 ( .A(n2211), .Y(n2212) );
  INVX1 U2295 ( .A(N120), .Y(n2213) );
  INVX4 U2296 ( .A(n2213), .Y(n2214) );
  INVX1 U2297 ( .A(N121), .Y(n2215) );
  INVX4 U2298 ( .A(n2215), .Y(n2216) );
  INVX1 U2299 ( .A(N122), .Y(n2217) );
  INVX4 U2300 ( .A(n2217), .Y(n2218) );
  INVX1 U2301 ( .A(N123), .Y(n2219) );
  INVX4 U2302 ( .A(n2219), .Y(n2220) );
  INVX1 U2303 ( .A(N124), .Y(n2221) );
  INVX4 U2304 ( .A(n2221), .Y(n2222) );
  INVX1 U2305 ( .A(N63), .Y(n2223) );
  INVX4 U2306 ( .A(n2223), .Y(n2224) );
  INVX1 U2307 ( .A(N94), .Y(n2225) );
  INVX4 U2308 ( .A(n2225), .Y(n2226) );
  INVX1 U2309 ( .A(N95), .Y(n2227) );
  INVX4 U2310 ( .A(n2227), .Y(n2228) );
  INVX1 U2311 ( .A(N96), .Y(n2229) );
  INVX4 U2312 ( .A(n2229), .Y(n2230) );
  INVX1 U2313 ( .A(N97), .Y(n2231) );
  INVX4 U2314 ( .A(n2231), .Y(n2232) );
  INVX1 U2315 ( .A(N98), .Y(n2233) );
  INVX4 U2316 ( .A(n2233), .Y(n2234) );
  INVX1 U2317 ( .A(N99), .Y(n2235) );
  INVX4 U2318 ( .A(n2235), .Y(n2236) );
  OR2X1 U2319 ( .A(address[7]), .B(address[6]), .Y(n2237) );
  AOI21X1 U2320 ( .A(address[5]), .B(address[4]), .C(n2237), .Y(N128) );
endmodule

